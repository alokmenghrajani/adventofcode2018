module delta_test;

  reg [25:0][7:0] a;
  reg [25:0][7:0] b;
  wire [5:0] r;

  delta dut (.a(a), .b(b), .r(r));

  initial begin
    $display("start");

    a[0] = 119; a[1] = 108; a[2] = 112; a[3] = 105; a[4] = 111; a[5] = 103; a[6] = 115; a[7] = 118; a[8] = 100; a[9] = 102; a[10] = 101; a[11] = 99; a[12] = 106; a[13] = 100; a[14] = 113; a[15] = 109; a[16] = 110; a[17] = 120; a[18] = 97; a[19] = 107; a[20] = 117; a[21] = 100; a[22] = 114; a[23] = 104; a[24] = 98; a[25] = 122;
    b[0] = 119; b[1] = 115; b[2] = 112; b[3] = 105; b[4] = 111; b[5] = 103; b[6] = 115; b[7] = 106; b[8] = 100; b[9] = 102; b[10] = 101; b[11] = 99; b[12] = 106; b[13] = 100; b[14] = 113; b[15] = 109; b[16] = 110; b[17] = 120; b[18] = 97; b[19] = 107; b[20] = 117; b[21] = 100; b[22] = 114; b[23] = 104; b[24] = 98; b[25] = 122; #10
    if (r != 24)
      $display("failed a=%b", a, ", b=%b", b, ", r=", r);

    $display("done");
  end

endmodule
