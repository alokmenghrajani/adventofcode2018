module field (
  input wire clk,
  input wire en,
  output wire [2499:0] trees,
  output wire [2499:0] lumberyards
);

acre acre_0_0 (.clk(clk), .en(en), .top_left(2'b0), .top(2'b0), .top_right(2'b0), .left(2'b0), .right({trees[1], lumberyards[1]}), .bottom_left(2'b0), .bottom({trees[50], lumberyards[50]}), .bottom_right({trees[51], lumberyards[51]}), .init(2'b00), .state({trees[0], lumberyards[0]}));
acre acre_0_1 (.clk(clk), .en(en), .top_left(2'b0), .top(2'b0), .top_right(2'b0), .left({trees[0], lumberyards[0]}), .right({trees[2], lumberyards[2]}), .bottom_left({trees[50], lumberyards[50]}), .bottom({trees[51], lumberyards[51]}), .bottom_right({trees[52], lumberyards[52]}), .init(2'b10), .state({trees[1], lumberyards[1]}));
acre acre_0_2 (.clk(clk), .en(en), .top_left(2'b0), .top(2'b0), .top_right(2'b0), .left({trees[1], lumberyards[1]}), .right({trees[3], lumberyards[3]}), .bottom_left({trees[51], lumberyards[51]}), .bottom({trees[52], lumberyards[52]}), .bottom_right({trees[53], lumberyards[53]}), .init(2'b00), .state({trees[2], lumberyards[2]}));
acre acre_0_3 (.clk(clk), .en(en), .top_left(2'b0), .top(2'b0), .top_right(2'b0), .left({trees[2], lumberyards[2]}), .right({trees[4], lumberyards[4]}), .bottom_left({trees[52], lumberyards[52]}), .bottom({trees[53], lumberyards[53]}), .bottom_right({trees[54], lumberyards[54]}), .init(2'b00), .state({trees[3], lumberyards[3]}));
acre acre_0_4 (.clk(clk), .en(en), .top_left(2'b0), .top(2'b0), .top_right(2'b0), .left({trees[3], lumberyards[3]}), .right({trees[5], lumberyards[5]}), .bottom_left({trees[53], lumberyards[53]}), .bottom({trees[54], lumberyards[54]}), .bottom_right({trees[55], lumberyards[55]}), .init(2'b00), .state({trees[4], lumberyards[4]}));
acre acre_0_5 (.clk(clk), .en(en), .top_left(2'b0), .top(2'b0), .top_right(2'b0), .left({trees[4], lumberyards[4]}), .right({trees[6], lumberyards[6]}), .bottom_left({trees[54], lumberyards[54]}), .bottom({trees[55], lumberyards[55]}), .bottom_right({trees[56], lumberyards[56]}), .init(2'b10), .state({trees[5], lumberyards[5]}));
acre acre_0_6 (.clk(clk), .en(en), .top_left(2'b0), .top(2'b0), .top_right(2'b0), .left({trees[5], lumberyards[5]}), .right({trees[7], lumberyards[7]}), .bottom_left({trees[55], lumberyards[55]}), .bottom({trees[56], lumberyards[56]}), .bottom_right({trees[57], lumberyards[57]}), .init(2'b00), .state({trees[6], lumberyards[6]}));
acre acre_0_7 (.clk(clk), .en(en), .top_left(2'b0), .top(2'b0), .top_right(2'b0), .left({trees[6], lumberyards[6]}), .right({trees[8], lumberyards[8]}), .bottom_left({trees[56], lumberyards[56]}), .bottom({trees[57], lumberyards[57]}), .bottom_right({trees[58], lumberyards[58]}), .init(2'b00), .state({trees[7], lumberyards[7]}));
acre acre_0_8 (.clk(clk), .en(en), .top_left(2'b0), .top(2'b0), .top_right(2'b0), .left({trees[7], lumberyards[7]}), .right({trees[9], lumberyards[9]}), .bottom_left({trees[57], lumberyards[57]}), .bottom({trees[58], lumberyards[58]}), .bottom_right({trees[59], lumberyards[59]}), .init(2'b10), .state({trees[8], lumberyards[8]}));
acre acre_0_9 (.clk(clk), .en(en), .top_left(2'b0), .top(2'b0), .top_right(2'b0), .left({trees[8], lumberyards[8]}), .right({trees[10], lumberyards[10]}), .bottom_left({trees[58], lumberyards[58]}), .bottom({trees[59], lumberyards[59]}), .bottom_right({trees[60], lumberyards[60]}), .init(2'b01), .state({trees[9], lumberyards[9]}));
acre acre_0_10 (.clk(clk), .en(en), .top_left(2'b0), .top(2'b0), .top_right(2'b0), .left({trees[9], lumberyards[9]}), .right({trees[11], lumberyards[11]}), .bottom_left({trees[59], lumberyards[59]}), .bottom({trees[60], lumberyards[60]}), .bottom_right({trees[61], lumberyards[61]}), .init(2'b01), .state({trees[10], lumberyards[10]}));
acre acre_0_11 (.clk(clk), .en(en), .top_left(2'b0), .top(2'b0), .top_right(2'b0), .left({trees[10], lumberyards[10]}), .right({trees[12], lumberyards[12]}), .bottom_left({trees[60], lumberyards[60]}), .bottom({trees[61], lumberyards[61]}), .bottom_right({trees[62], lumberyards[62]}), .init(2'b00), .state({trees[11], lumberyards[11]}));
acre acre_0_12 (.clk(clk), .en(en), .top_left(2'b0), .top(2'b0), .top_right(2'b0), .left({trees[11], lumberyards[11]}), .right({trees[13], lumberyards[13]}), .bottom_left({trees[61], lumberyards[61]}), .bottom({trees[62], lumberyards[62]}), .bottom_right({trees[63], lumberyards[63]}), .init(2'b01), .state({trees[12], lumberyards[12]}));
acre acre_0_13 (.clk(clk), .en(en), .top_left(2'b0), .top(2'b0), .top_right(2'b0), .left({trees[12], lumberyards[12]}), .right({trees[14], lumberyards[14]}), .bottom_left({trees[62], lumberyards[62]}), .bottom({trees[63], lumberyards[63]}), .bottom_right({trees[64], lumberyards[64]}), .init(2'b00), .state({trees[13], lumberyards[13]}));
acre acre_0_14 (.clk(clk), .en(en), .top_left(2'b0), .top(2'b0), .top_right(2'b0), .left({trees[13], lumberyards[13]}), .right({trees[15], lumberyards[15]}), .bottom_left({trees[63], lumberyards[63]}), .bottom({trees[64], lumberyards[64]}), .bottom_right({trees[65], lumberyards[65]}), .init(2'b10), .state({trees[14], lumberyards[14]}));
acre acre_0_15 (.clk(clk), .en(en), .top_left(2'b0), .top(2'b0), .top_right(2'b0), .left({trees[14], lumberyards[14]}), .right({trees[16], lumberyards[16]}), .bottom_left({trees[64], lumberyards[64]}), .bottom({trees[65], lumberyards[65]}), .bottom_right({trees[66], lumberyards[66]}), .init(2'b01), .state({trees[15], lumberyards[15]}));
acre acre_0_16 (.clk(clk), .en(en), .top_left(2'b0), .top(2'b0), .top_right(2'b0), .left({trees[15], lumberyards[15]}), .right({trees[17], lumberyards[17]}), .bottom_left({trees[65], lumberyards[65]}), .bottom({trees[66], lumberyards[66]}), .bottom_right({trees[67], lumberyards[67]}), .init(2'b01), .state({trees[16], lumberyards[16]}));
acre acre_0_17 (.clk(clk), .en(en), .top_left(2'b0), .top(2'b0), .top_right(2'b0), .left({trees[16], lumberyards[16]}), .right({trees[18], lumberyards[18]}), .bottom_left({trees[66], lumberyards[66]}), .bottom({trees[67], lumberyards[67]}), .bottom_right({trees[68], lumberyards[68]}), .init(2'b00), .state({trees[17], lumberyards[17]}));
acre acre_0_18 (.clk(clk), .en(en), .top_left(2'b0), .top(2'b0), .top_right(2'b0), .left({trees[17], lumberyards[17]}), .right({trees[19], lumberyards[19]}), .bottom_left({trees[67], lumberyards[67]}), .bottom({trees[68], lumberyards[68]}), .bottom_right({trees[69], lumberyards[69]}), .init(2'b00), .state({trees[18], lumberyards[18]}));
acre acre_0_19 (.clk(clk), .en(en), .top_left(2'b0), .top(2'b0), .top_right(2'b0), .left({trees[18], lumberyards[18]}), .right({trees[20], lumberyards[20]}), .bottom_left({trees[68], lumberyards[68]}), .bottom({trees[69], lumberyards[69]}), .bottom_right({trees[70], lumberyards[70]}), .init(2'b00), .state({trees[19], lumberyards[19]}));
acre acre_0_20 (.clk(clk), .en(en), .top_left(2'b0), .top(2'b0), .top_right(2'b0), .left({trees[19], lumberyards[19]}), .right({trees[21], lumberyards[21]}), .bottom_left({trees[69], lumberyards[69]}), .bottom({trees[70], lumberyards[70]}), .bottom_right({trees[71], lumberyards[71]}), .init(2'b01), .state({trees[20], lumberyards[20]}));
acre acre_0_21 (.clk(clk), .en(en), .top_left(2'b0), .top(2'b0), .top_right(2'b0), .left({trees[20], lumberyards[20]}), .right({trees[22], lumberyards[22]}), .bottom_left({trees[70], lumberyards[70]}), .bottom({trees[71], lumberyards[71]}), .bottom_right({trees[72], lumberyards[72]}), .init(2'b00), .state({trees[21], lumberyards[21]}));
acre acre_0_22 (.clk(clk), .en(en), .top_left(2'b0), .top(2'b0), .top_right(2'b0), .left({trees[21], lumberyards[21]}), .right({trees[23], lumberyards[23]}), .bottom_left({trees[71], lumberyards[71]}), .bottom({trees[72], lumberyards[72]}), .bottom_right({trees[73], lumberyards[73]}), .init(2'b10), .state({trees[22], lumberyards[22]}));
acre acre_0_23 (.clk(clk), .en(en), .top_left(2'b0), .top(2'b0), .top_right(2'b0), .left({trees[22], lumberyards[22]}), .right({trees[24], lumberyards[24]}), .bottom_left({trees[72], lumberyards[72]}), .bottom({trees[73], lumberyards[73]}), .bottom_right({trees[74], lumberyards[74]}), .init(2'b00), .state({trees[23], lumberyards[23]}));
acre acre_0_24 (.clk(clk), .en(en), .top_left(2'b0), .top(2'b0), .top_right(2'b0), .left({trees[23], lumberyards[23]}), .right({trees[25], lumberyards[25]}), .bottom_left({trees[73], lumberyards[73]}), .bottom({trees[74], lumberyards[74]}), .bottom_right({trees[75], lumberyards[75]}), .init(2'b00), .state({trees[24], lumberyards[24]}));
acre acre_0_25 (.clk(clk), .en(en), .top_left(2'b0), .top(2'b0), .top_right(2'b0), .left({trees[24], lumberyards[24]}), .right({trees[26], lumberyards[26]}), .bottom_left({trees[74], lumberyards[74]}), .bottom({trees[75], lumberyards[75]}), .bottom_right({trees[76], lumberyards[76]}), .init(2'b00), .state({trees[25], lumberyards[25]}));
acre acre_0_26 (.clk(clk), .en(en), .top_left(2'b0), .top(2'b0), .top_right(2'b0), .left({trees[25], lumberyards[25]}), .right({trees[27], lumberyards[27]}), .bottom_left({trees[75], lumberyards[75]}), .bottom({trees[76], lumberyards[76]}), .bottom_right({trees[77], lumberyards[77]}), .init(2'b00), .state({trees[26], lumberyards[26]}));
acre acre_0_27 (.clk(clk), .en(en), .top_left(2'b0), .top(2'b0), .top_right(2'b0), .left({trees[26], lumberyards[26]}), .right({trees[28], lumberyards[28]}), .bottom_left({trees[76], lumberyards[76]}), .bottom({trees[77], lumberyards[77]}), .bottom_right({trees[78], lumberyards[78]}), .init(2'b00), .state({trees[27], lumberyards[27]}));
acre acre_0_28 (.clk(clk), .en(en), .top_left(2'b0), .top(2'b0), .top_right(2'b0), .left({trees[27], lumberyards[27]}), .right({trees[29], lumberyards[29]}), .bottom_left({trees[77], lumberyards[77]}), .bottom({trees[78], lumberyards[78]}), .bottom_right({trees[79], lumberyards[79]}), .init(2'b00), .state({trees[28], lumberyards[28]}));
acre acre_0_29 (.clk(clk), .en(en), .top_left(2'b0), .top(2'b0), .top_right(2'b0), .left({trees[28], lumberyards[28]}), .right({trees[30], lumberyards[30]}), .bottom_left({trees[78], lumberyards[78]}), .bottom({trees[79], lumberyards[79]}), .bottom_right({trees[80], lumberyards[80]}), .init(2'b00), .state({trees[29], lumberyards[29]}));
acre acre_0_30 (.clk(clk), .en(en), .top_left(2'b0), .top(2'b0), .top_right(2'b0), .left({trees[29], lumberyards[29]}), .right({trees[31], lumberyards[31]}), .bottom_left({trees[79], lumberyards[79]}), .bottom({trees[80], lumberyards[80]}), .bottom_right({trees[81], lumberyards[81]}), .init(2'b00), .state({trees[30], lumberyards[30]}));
acre acre_0_31 (.clk(clk), .en(en), .top_left(2'b0), .top(2'b0), .top_right(2'b0), .left({trees[30], lumberyards[30]}), .right({trees[32], lumberyards[32]}), .bottom_left({trees[80], lumberyards[80]}), .bottom({trees[81], lumberyards[81]}), .bottom_right({trees[82], lumberyards[82]}), .init(2'b10), .state({trees[31], lumberyards[31]}));
acre acre_0_32 (.clk(clk), .en(en), .top_left(2'b0), .top(2'b0), .top_right(2'b0), .left({trees[31], lumberyards[31]}), .right({trees[33], lumberyards[33]}), .bottom_left({trees[81], lumberyards[81]}), .bottom({trees[82], lumberyards[82]}), .bottom_right({trees[83], lumberyards[83]}), .init(2'b00), .state({trees[32], lumberyards[32]}));
acre acre_0_33 (.clk(clk), .en(en), .top_left(2'b0), .top(2'b0), .top_right(2'b0), .left({trees[32], lumberyards[32]}), .right({trees[34], lumberyards[34]}), .bottom_left({trees[82], lumberyards[82]}), .bottom({trees[83], lumberyards[83]}), .bottom_right({trees[84], lumberyards[84]}), .init(2'b00), .state({trees[33], lumberyards[33]}));
acre acre_0_34 (.clk(clk), .en(en), .top_left(2'b0), .top(2'b0), .top_right(2'b0), .left({trees[33], lumberyards[33]}), .right({trees[35], lumberyards[35]}), .bottom_left({trees[83], lumberyards[83]}), .bottom({trees[84], lumberyards[84]}), .bottom_right({trees[85], lumberyards[85]}), .init(2'b10), .state({trees[34], lumberyards[34]}));
acre acre_0_35 (.clk(clk), .en(en), .top_left(2'b0), .top(2'b0), .top_right(2'b0), .left({trees[34], lumberyards[34]}), .right({trees[36], lumberyards[36]}), .bottom_left({trees[84], lumberyards[84]}), .bottom({trees[85], lumberyards[85]}), .bottom_right({trees[86], lumberyards[86]}), .init(2'b00), .state({trees[35], lumberyards[35]}));
acre acre_0_36 (.clk(clk), .en(en), .top_left(2'b0), .top(2'b0), .top_right(2'b0), .left({trees[35], lumberyards[35]}), .right({trees[37], lumberyards[37]}), .bottom_left({trees[85], lumberyards[85]}), .bottom({trees[86], lumberyards[86]}), .bottom_right({trees[87], lumberyards[87]}), .init(2'b00), .state({trees[36], lumberyards[36]}));
acre acre_0_37 (.clk(clk), .en(en), .top_left(2'b0), .top(2'b0), .top_right(2'b0), .left({trees[36], lumberyards[36]}), .right({trees[38], lumberyards[38]}), .bottom_left({trees[86], lumberyards[86]}), .bottom({trees[87], lumberyards[87]}), .bottom_right({trees[88], lumberyards[88]}), .init(2'b00), .state({trees[37], lumberyards[37]}));
acre acre_0_38 (.clk(clk), .en(en), .top_left(2'b0), .top(2'b0), .top_right(2'b0), .left({trees[37], lumberyards[37]}), .right({trees[39], lumberyards[39]}), .bottom_left({trees[87], lumberyards[87]}), .bottom({trees[88], lumberyards[88]}), .bottom_right({trees[89], lumberyards[89]}), .init(2'b01), .state({trees[38], lumberyards[38]}));
acre acre_0_39 (.clk(clk), .en(en), .top_left(2'b0), .top(2'b0), .top_right(2'b0), .left({trees[38], lumberyards[38]}), .right({trees[40], lumberyards[40]}), .bottom_left({trees[88], lumberyards[88]}), .bottom({trees[89], lumberyards[89]}), .bottom_right({trees[90], lumberyards[90]}), .init(2'b00), .state({trees[39], lumberyards[39]}));
acre acre_0_40 (.clk(clk), .en(en), .top_left(2'b0), .top(2'b0), .top_right(2'b0), .left({trees[39], lumberyards[39]}), .right({trees[41], lumberyards[41]}), .bottom_left({trees[89], lumberyards[89]}), .bottom({trees[90], lumberyards[90]}), .bottom_right({trees[91], lumberyards[91]}), .init(2'b00), .state({trees[40], lumberyards[40]}));
acre acre_0_41 (.clk(clk), .en(en), .top_left(2'b0), .top(2'b0), .top_right(2'b0), .left({trees[40], lumberyards[40]}), .right({trees[42], lumberyards[42]}), .bottom_left({trees[90], lumberyards[90]}), .bottom({trees[91], lumberyards[91]}), .bottom_right({trees[92], lumberyards[92]}), .init(2'b10), .state({trees[41], lumberyards[41]}));
acre acre_0_42 (.clk(clk), .en(en), .top_left(2'b0), .top(2'b0), .top_right(2'b0), .left({trees[41], lumberyards[41]}), .right({trees[43], lumberyards[43]}), .bottom_left({trees[91], lumberyards[91]}), .bottom({trees[92], lumberyards[92]}), .bottom_right({trees[93], lumberyards[93]}), .init(2'b01), .state({trees[42], lumberyards[42]}));
acre acre_0_43 (.clk(clk), .en(en), .top_left(2'b0), .top(2'b0), .top_right(2'b0), .left({trees[42], lumberyards[42]}), .right({trees[44], lumberyards[44]}), .bottom_left({trees[92], lumberyards[92]}), .bottom({trees[93], lumberyards[93]}), .bottom_right({trees[94], lumberyards[94]}), .init(2'b01), .state({trees[43], lumberyards[43]}));
acre acre_0_44 (.clk(clk), .en(en), .top_left(2'b0), .top(2'b0), .top_right(2'b0), .left({trees[43], lumberyards[43]}), .right({trees[45], lumberyards[45]}), .bottom_left({trees[93], lumberyards[93]}), .bottom({trees[94], lumberyards[94]}), .bottom_right({trees[95], lumberyards[95]}), .init(2'b00), .state({trees[44], lumberyards[44]}));
acre acre_0_45 (.clk(clk), .en(en), .top_left(2'b0), .top(2'b0), .top_right(2'b0), .left({trees[44], lumberyards[44]}), .right({trees[46], lumberyards[46]}), .bottom_left({trees[94], lumberyards[94]}), .bottom({trees[95], lumberyards[95]}), .bottom_right({trees[96], lumberyards[96]}), .init(2'b10), .state({trees[45], lumberyards[45]}));
acre acre_0_46 (.clk(clk), .en(en), .top_left(2'b0), .top(2'b0), .top_right(2'b0), .left({trees[45], lumberyards[45]}), .right({trees[47], lumberyards[47]}), .bottom_left({trees[95], lumberyards[95]}), .bottom({trees[96], lumberyards[96]}), .bottom_right({trees[97], lumberyards[97]}), .init(2'b00), .state({trees[46], lumberyards[46]}));
acre acre_0_47 (.clk(clk), .en(en), .top_left(2'b0), .top(2'b0), .top_right(2'b0), .left({trees[46], lumberyards[46]}), .right({trees[48], lumberyards[48]}), .bottom_left({trees[96], lumberyards[96]}), .bottom({trees[97], lumberyards[97]}), .bottom_right({trees[98], lumberyards[98]}), .init(2'b00), .state({trees[47], lumberyards[47]}));
acre acre_0_48 (.clk(clk), .en(en), .top_left(2'b0), .top(2'b0), .top_right(2'b0), .left({trees[47], lumberyards[47]}), .right({trees[49], lumberyards[49]}), .bottom_left({trees[97], lumberyards[97]}), .bottom({trees[98], lumberyards[98]}), .bottom_right({trees[99], lumberyards[99]}), .init(2'b00), .state({trees[48], lumberyards[48]}));
acre acre_0_49 (.clk(clk), .en(en), .top_left(2'b0), .top(2'b0), .top_right(2'b0), .left({trees[48], lumberyards[48]}), .right(2'b0), .bottom_left({trees[98], lumberyards[98]}), .bottom({trees[99], lumberyards[99]}), .bottom_right(2'b0), .init(2'b00), .state({trees[49], lumberyards[49]}));
acre acre_1_0 (.clk(clk), .en(en), .top_left(2'b0), .top({trees[0], lumberyards[0]}), .top_right({trees[1], lumberyards[1]}), .left(2'b0), .right({trees[51], lumberyards[51]}), .bottom_left(2'b0), .bottom({trees[100], lumberyards[100]}), .bottom_right({trees[101], lumberyards[101]}), .init(2'b00), .state({trees[50], lumberyards[50]}));
acre acre_1_1 (.clk(clk), .en(en), .top_left({trees[0], lumberyards[0]}), .top({trees[1], lumberyards[1]}), .top_right({trees[2], lumberyards[2]}), .left({trees[50], lumberyards[50]}), .right({trees[52], lumberyards[52]}), .bottom_left({trees[100], lumberyards[100]}), .bottom({trees[101], lumberyards[101]}), .bottom_right({trees[102], lumberyards[102]}), .init(2'b00), .state({trees[51], lumberyards[51]}));
acre acre_1_2 (.clk(clk), .en(en), .top_left({trees[1], lumberyards[1]}), .top({trees[2], lumberyards[2]}), .top_right({trees[3], lumberyards[3]}), .left({trees[51], lumberyards[51]}), .right({trees[53], lumberyards[53]}), .bottom_left({trees[101], lumberyards[101]}), .bottom({trees[102], lumberyards[102]}), .bottom_right({trees[103], lumberyards[103]}), .init(2'b01), .state({trees[52], lumberyards[52]}));
acre acre_1_3 (.clk(clk), .en(en), .top_left({trees[2], lumberyards[2]}), .top({trees[3], lumberyards[3]}), .top_right({trees[4], lumberyards[4]}), .left({trees[52], lumberyards[52]}), .right({trees[54], lumberyards[54]}), .bottom_left({trees[102], lumberyards[102]}), .bottom({trees[103], lumberyards[103]}), .bottom_right({trees[104], lumberyards[104]}), .init(2'b00), .state({trees[53], lumberyards[53]}));
acre acre_1_4 (.clk(clk), .en(en), .top_left({trees[3], lumberyards[3]}), .top({trees[4], lumberyards[4]}), .top_right({trees[5], lumberyards[5]}), .left({trees[53], lumberyards[53]}), .right({trees[55], lumberyards[55]}), .bottom_left({trees[103], lumberyards[103]}), .bottom({trees[104], lumberyards[104]}), .bottom_right({trees[105], lumberyards[105]}), .init(2'b00), .state({trees[54], lumberyards[54]}));
acre acre_1_5 (.clk(clk), .en(en), .top_left({trees[4], lumberyards[4]}), .top({trees[5], lumberyards[5]}), .top_right({trees[6], lumberyards[6]}), .left({trees[54], lumberyards[54]}), .right({trees[56], lumberyards[56]}), .bottom_left({trees[104], lumberyards[104]}), .bottom({trees[105], lumberyards[105]}), .bottom_right({trees[106], lumberyards[106]}), .init(2'b00), .state({trees[55], lumberyards[55]}));
acre acre_1_6 (.clk(clk), .en(en), .top_left({trees[5], lumberyards[5]}), .top({trees[6], lumberyards[6]}), .top_right({trees[7], lumberyards[7]}), .left({trees[55], lumberyards[55]}), .right({trees[57], lumberyards[57]}), .bottom_left({trees[105], lumberyards[105]}), .bottom({trees[106], lumberyards[106]}), .bottom_right({trees[107], lumberyards[107]}), .init(2'b00), .state({trees[56], lumberyards[56]}));
acre acre_1_7 (.clk(clk), .en(en), .top_left({trees[6], lumberyards[6]}), .top({trees[7], lumberyards[7]}), .top_right({trees[8], lumberyards[8]}), .left({trees[56], lumberyards[56]}), .right({trees[58], lumberyards[58]}), .bottom_left({trees[106], lumberyards[106]}), .bottom({trees[107], lumberyards[107]}), .bottom_right({trees[108], lumberyards[108]}), .init(2'b01), .state({trees[57], lumberyards[57]}));
acre acre_1_8 (.clk(clk), .en(en), .top_left({trees[7], lumberyards[7]}), .top({trees[8], lumberyards[8]}), .top_right({trees[9], lumberyards[9]}), .left({trees[57], lumberyards[57]}), .right({trees[59], lumberyards[59]}), .bottom_left({trees[107], lumberyards[107]}), .bottom({trees[108], lumberyards[108]}), .bottom_right({trees[109], lumberyards[109]}), .init(2'b00), .state({trees[58], lumberyards[58]}));
acre acre_1_9 (.clk(clk), .en(en), .top_left({trees[8], lumberyards[8]}), .top({trees[9], lumberyards[9]}), .top_right({trees[10], lumberyards[10]}), .left({trees[58], lumberyards[58]}), .right({trees[60], lumberyards[60]}), .bottom_left({trees[108], lumberyards[108]}), .bottom({trees[109], lumberyards[109]}), .bottom_right({trees[110], lumberyards[110]}), .init(2'b10), .state({trees[59], lumberyards[59]}));
acre acre_1_10 (.clk(clk), .en(en), .top_left({trees[9], lumberyards[9]}), .top({trees[10], lumberyards[10]}), .top_right({trees[11], lumberyards[11]}), .left({trees[59], lumberyards[59]}), .right({trees[61], lumberyards[61]}), .bottom_left({trees[109], lumberyards[109]}), .bottom({trees[110], lumberyards[110]}), .bottom_right({trees[111], lumberyards[111]}), .init(2'b00), .state({trees[60], lumberyards[60]}));
acre acre_1_11 (.clk(clk), .en(en), .top_left({trees[10], lumberyards[10]}), .top({trees[11], lumberyards[11]}), .top_right({trees[12], lumberyards[12]}), .left({trees[60], lumberyards[60]}), .right({trees[62], lumberyards[62]}), .bottom_left({trees[110], lumberyards[110]}), .bottom({trees[111], lumberyards[111]}), .bottom_right({trees[112], lumberyards[112]}), .init(2'b00), .state({trees[61], lumberyards[61]}));
acre acre_1_12 (.clk(clk), .en(en), .top_left({trees[11], lumberyards[11]}), .top({trees[12], lumberyards[12]}), .top_right({trees[13], lumberyards[13]}), .left({trees[61], lumberyards[61]}), .right({trees[63], lumberyards[63]}), .bottom_left({trees[111], lumberyards[111]}), .bottom({trees[112], lumberyards[112]}), .bottom_right({trees[113], lumberyards[113]}), .init(2'b00), .state({trees[62], lumberyards[62]}));
acre acre_1_13 (.clk(clk), .en(en), .top_left({trees[12], lumberyards[12]}), .top({trees[13], lumberyards[13]}), .top_right({trees[14], lumberyards[14]}), .left({trees[62], lumberyards[62]}), .right({trees[64], lumberyards[64]}), .bottom_left({trees[112], lumberyards[112]}), .bottom({trees[113], lumberyards[113]}), .bottom_right({trees[114], lumberyards[114]}), .init(2'b00), .state({trees[63], lumberyards[63]}));
acre acre_1_14 (.clk(clk), .en(en), .top_left({trees[13], lumberyards[13]}), .top({trees[14], lumberyards[14]}), .top_right({trees[15], lumberyards[15]}), .left({trees[63], lumberyards[63]}), .right({trees[65], lumberyards[65]}), .bottom_left({trees[113], lumberyards[113]}), .bottom({trees[114], lumberyards[114]}), .bottom_right({trees[115], lumberyards[115]}), .init(2'b00), .state({trees[64], lumberyards[64]}));
acre acre_1_15 (.clk(clk), .en(en), .top_left({trees[14], lumberyards[14]}), .top({trees[15], lumberyards[15]}), .top_right({trees[16], lumberyards[16]}), .left({trees[64], lumberyards[64]}), .right({trees[66], lumberyards[66]}), .bottom_left({trees[114], lumberyards[114]}), .bottom({trees[115], lumberyards[115]}), .bottom_right({trees[116], lumberyards[116]}), .init(2'b00), .state({trees[65], lumberyards[65]}));
acre acre_1_16 (.clk(clk), .en(en), .top_left({trees[15], lumberyards[15]}), .top({trees[16], lumberyards[16]}), .top_right({trees[17], lumberyards[17]}), .left({trees[65], lumberyards[65]}), .right({trees[67], lumberyards[67]}), .bottom_left({trees[115], lumberyards[115]}), .bottom({trees[116], lumberyards[116]}), .bottom_right({trees[117], lumberyards[117]}), .init(2'b00), .state({trees[66], lumberyards[66]}));
acre acre_1_17 (.clk(clk), .en(en), .top_left({trees[16], lumberyards[16]}), .top({trees[17], lumberyards[17]}), .top_right({trees[18], lumberyards[18]}), .left({trees[66], lumberyards[66]}), .right({trees[68], lumberyards[68]}), .bottom_left({trees[116], lumberyards[116]}), .bottom({trees[117], lumberyards[117]}), .bottom_right({trees[118], lumberyards[118]}), .init(2'b00), .state({trees[67], lumberyards[67]}));
acre acre_1_18 (.clk(clk), .en(en), .top_left({trees[17], lumberyards[17]}), .top({trees[18], lumberyards[18]}), .top_right({trees[19], lumberyards[19]}), .left({trees[67], lumberyards[67]}), .right({trees[69], lumberyards[69]}), .bottom_left({trees[117], lumberyards[117]}), .bottom({trees[118], lumberyards[118]}), .bottom_right({trees[119], lumberyards[119]}), .init(2'b00), .state({trees[68], lumberyards[68]}));
acre acre_1_19 (.clk(clk), .en(en), .top_left({trees[18], lumberyards[18]}), .top({trees[19], lumberyards[19]}), .top_right({trees[20], lumberyards[20]}), .left({trees[68], lumberyards[68]}), .right({trees[70], lumberyards[70]}), .bottom_left({trees[118], lumberyards[118]}), .bottom({trees[119], lumberyards[119]}), .bottom_right({trees[120], lumberyards[120]}), .init(2'b00), .state({trees[69], lumberyards[69]}));
acre acre_1_20 (.clk(clk), .en(en), .top_left({trees[19], lumberyards[19]}), .top({trees[20], lumberyards[20]}), .top_right({trees[21], lumberyards[21]}), .left({trees[69], lumberyards[69]}), .right({trees[71], lumberyards[71]}), .bottom_left({trees[119], lumberyards[119]}), .bottom({trees[120], lumberyards[120]}), .bottom_right({trees[121], lumberyards[121]}), .init(2'b10), .state({trees[70], lumberyards[70]}));
acre acre_1_21 (.clk(clk), .en(en), .top_left({trees[20], lumberyards[20]}), .top({trees[21], lumberyards[21]}), .top_right({trees[22], lumberyards[22]}), .left({trees[70], lumberyards[70]}), .right({trees[72], lumberyards[72]}), .bottom_left({trees[120], lumberyards[120]}), .bottom({trees[121], lumberyards[121]}), .bottom_right({trees[122], lumberyards[122]}), .init(2'b01), .state({trees[71], lumberyards[71]}));
acre acre_1_22 (.clk(clk), .en(en), .top_left({trees[21], lumberyards[21]}), .top({trees[22], lumberyards[22]}), .top_right({trees[23], lumberyards[23]}), .left({trees[71], lumberyards[71]}), .right({trees[73], lumberyards[73]}), .bottom_left({trees[121], lumberyards[121]}), .bottom({trees[122], lumberyards[122]}), .bottom_right({trees[123], lumberyards[123]}), .init(2'b00), .state({trees[72], lumberyards[72]}));
acre acre_1_23 (.clk(clk), .en(en), .top_left({trees[22], lumberyards[22]}), .top({trees[23], lumberyards[23]}), .top_right({trees[24], lumberyards[24]}), .left({trees[72], lumberyards[72]}), .right({trees[74], lumberyards[74]}), .bottom_left({trees[122], lumberyards[122]}), .bottom({trees[123], lumberyards[123]}), .bottom_right({trees[124], lumberyards[124]}), .init(2'b00), .state({trees[73], lumberyards[73]}));
acre acre_1_24 (.clk(clk), .en(en), .top_left({trees[23], lumberyards[23]}), .top({trees[24], lumberyards[24]}), .top_right({trees[25], lumberyards[25]}), .left({trees[73], lumberyards[73]}), .right({trees[75], lumberyards[75]}), .bottom_left({trees[123], lumberyards[123]}), .bottom({trees[124], lumberyards[124]}), .bottom_right({trees[125], lumberyards[125]}), .init(2'b00), .state({trees[74], lumberyards[74]}));
acre acre_1_25 (.clk(clk), .en(en), .top_left({trees[24], lumberyards[24]}), .top({trees[25], lumberyards[25]}), .top_right({trees[26], lumberyards[26]}), .left({trees[74], lumberyards[74]}), .right({trees[76], lumberyards[76]}), .bottom_left({trees[124], lumberyards[124]}), .bottom({trees[125], lumberyards[125]}), .bottom_right({trees[126], lumberyards[126]}), .init(2'b00), .state({trees[75], lumberyards[75]}));
acre acre_1_26 (.clk(clk), .en(en), .top_left({trees[25], lumberyards[25]}), .top({trees[26], lumberyards[26]}), .top_right({trees[27], lumberyards[27]}), .left({trees[75], lumberyards[75]}), .right({trees[77], lumberyards[77]}), .bottom_left({trees[125], lumberyards[125]}), .bottom({trees[126], lumberyards[126]}), .bottom_right({trees[127], lumberyards[127]}), .init(2'b00), .state({trees[76], lumberyards[76]}));
acre acre_1_27 (.clk(clk), .en(en), .top_left({trees[26], lumberyards[26]}), .top({trees[27], lumberyards[27]}), .top_right({trees[28], lumberyards[28]}), .left({trees[76], lumberyards[76]}), .right({trees[78], lumberyards[78]}), .bottom_left({trees[126], lumberyards[126]}), .bottom({trees[127], lumberyards[127]}), .bottom_right({trees[128], lumberyards[128]}), .init(2'b01), .state({trees[77], lumberyards[77]}));
acre acre_1_28 (.clk(clk), .en(en), .top_left({trees[27], lumberyards[27]}), .top({trees[28], lumberyards[28]}), .top_right({trees[29], lumberyards[29]}), .left({trees[77], lumberyards[77]}), .right({trees[79], lumberyards[79]}), .bottom_left({trees[127], lumberyards[127]}), .bottom({trees[128], lumberyards[128]}), .bottom_right({trees[129], lumberyards[129]}), .init(2'b01), .state({trees[78], lumberyards[78]}));
acre acre_1_29 (.clk(clk), .en(en), .top_left({trees[28], lumberyards[28]}), .top({trees[29], lumberyards[29]}), .top_right({trees[30], lumberyards[30]}), .left({trees[78], lumberyards[78]}), .right({trees[80], lumberyards[80]}), .bottom_left({trees[128], lumberyards[128]}), .bottom({trees[129], lumberyards[129]}), .bottom_right({trees[130], lumberyards[130]}), .init(2'b00), .state({trees[79], lumberyards[79]}));
acre acre_1_30 (.clk(clk), .en(en), .top_left({trees[29], lumberyards[29]}), .top({trees[30], lumberyards[30]}), .top_right({trees[31], lumberyards[31]}), .left({trees[79], lumberyards[79]}), .right({trees[81], lumberyards[81]}), .bottom_left({trees[129], lumberyards[129]}), .bottom({trees[130], lumberyards[130]}), .bottom_right({trees[131], lumberyards[131]}), .init(2'b00), .state({trees[80], lumberyards[80]}));
acre acre_1_31 (.clk(clk), .en(en), .top_left({trees[30], lumberyards[30]}), .top({trees[31], lumberyards[31]}), .top_right({trees[32], lumberyards[32]}), .left({trees[80], lumberyards[80]}), .right({trees[82], lumberyards[82]}), .bottom_left({trees[130], lumberyards[130]}), .bottom({trees[131], lumberyards[131]}), .bottom_right({trees[132], lumberyards[132]}), .init(2'b10), .state({trees[81], lumberyards[81]}));
acre acre_1_32 (.clk(clk), .en(en), .top_left({trees[31], lumberyards[31]}), .top({trees[32], lumberyards[32]}), .top_right({trees[33], lumberyards[33]}), .left({trees[81], lumberyards[81]}), .right({trees[83], lumberyards[83]}), .bottom_left({trees[131], lumberyards[131]}), .bottom({trees[132], lumberyards[132]}), .bottom_right({trees[133], lumberyards[133]}), .init(2'b00), .state({trees[82], lumberyards[82]}));
acre acre_1_33 (.clk(clk), .en(en), .top_left({trees[32], lumberyards[32]}), .top({trees[33], lumberyards[33]}), .top_right({trees[34], lumberyards[34]}), .left({trees[82], lumberyards[82]}), .right({trees[84], lumberyards[84]}), .bottom_left({trees[132], lumberyards[132]}), .bottom({trees[133], lumberyards[133]}), .bottom_right({trees[134], lumberyards[134]}), .init(2'b00), .state({trees[83], lumberyards[83]}));
acre acre_1_34 (.clk(clk), .en(en), .top_left({trees[33], lumberyards[33]}), .top({trees[34], lumberyards[34]}), .top_right({trees[35], lumberyards[35]}), .left({trees[83], lumberyards[83]}), .right({trees[85], lumberyards[85]}), .bottom_left({trees[133], lumberyards[133]}), .bottom({trees[134], lumberyards[134]}), .bottom_right({trees[135], lumberyards[135]}), .init(2'b00), .state({trees[84], lumberyards[84]}));
acre acre_1_35 (.clk(clk), .en(en), .top_left({trees[34], lumberyards[34]}), .top({trees[35], lumberyards[35]}), .top_right({trees[36], lumberyards[36]}), .left({trees[84], lumberyards[84]}), .right({trees[86], lumberyards[86]}), .bottom_left({trees[134], lumberyards[134]}), .bottom({trees[135], lumberyards[135]}), .bottom_right({trees[136], lumberyards[136]}), .init(2'b10), .state({trees[85], lumberyards[85]}));
acre acre_1_36 (.clk(clk), .en(en), .top_left({trees[35], lumberyards[35]}), .top({trees[36], lumberyards[36]}), .top_right({trees[37], lumberyards[37]}), .left({trees[85], lumberyards[85]}), .right({trees[87], lumberyards[87]}), .bottom_left({trees[135], lumberyards[135]}), .bottom({trees[136], lumberyards[136]}), .bottom_right({trees[137], lumberyards[137]}), .init(2'b01), .state({trees[86], lumberyards[86]}));
acre acre_1_37 (.clk(clk), .en(en), .top_left({trees[36], lumberyards[36]}), .top({trees[37], lumberyards[37]}), .top_right({trees[38], lumberyards[38]}), .left({trees[86], lumberyards[86]}), .right({trees[88], lumberyards[88]}), .bottom_left({trees[136], lumberyards[136]}), .bottom({trees[137], lumberyards[137]}), .bottom_right({trees[138], lumberyards[138]}), .init(2'b10), .state({trees[87], lumberyards[87]}));
acre acre_1_38 (.clk(clk), .en(en), .top_left({trees[37], lumberyards[37]}), .top({trees[38], lumberyards[38]}), .top_right({trees[39], lumberyards[39]}), .left({trees[87], lumberyards[87]}), .right({trees[89], lumberyards[89]}), .bottom_left({trees[137], lumberyards[137]}), .bottom({trees[138], lumberyards[138]}), .bottom_right({trees[139], lumberyards[139]}), .init(2'b10), .state({trees[88], lumberyards[88]}));
acre acre_1_39 (.clk(clk), .en(en), .top_left({trees[38], lumberyards[38]}), .top({trees[39], lumberyards[39]}), .top_right({trees[40], lumberyards[40]}), .left({trees[88], lumberyards[88]}), .right({trees[90], lumberyards[90]}), .bottom_left({trees[138], lumberyards[138]}), .bottom({trees[139], lumberyards[139]}), .bottom_right({trees[140], lumberyards[140]}), .init(2'b00), .state({trees[89], lumberyards[89]}));
acre acre_1_40 (.clk(clk), .en(en), .top_left({trees[39], lumberyards[39]}), .top({trees[40], lumberyards[40]}), .top_right({trees[41], lumberyards[41]}), .left({trees[89], lumberyards[89]}), .right({trees[91], lumberyards[91]}), .bottom_left({trees[139], lumberyards[139]}), .bottom({trees[140], lumberyards[140]}), .bottom_right({trees[141], lumberyards[141]}), .init(2'b00), .state({trees[90], lumberyards[90]}));
acre acre_1_41 (.clk(clk), .en(en), .top_left({trees[40], lumberyards[40]}), .top({trees[41], lumberyards[41]}), .top_right({trees[42], lumberyards[42]}), .left({trees[90], lumberyards[90]}), .right({trees[92], lumberyards[92]}), .bottom_left({trees[140], lumberyards[140]}), .bottom({trees[141], lumberyards[141]}), .bottom_right({trees[142], lumberyards[142]}), .init(2'b00), .state({trees[91], lumberyards[91]}));
acre acre_1_42 (.clk(clk), .en(en), .top_left({trees[41], lumberyards[41]}), .top({trees[42], lumberyards[42]}), .top_right({trees[43], lumberyards[43]}), .left({trees[91], lumberyards[91]}), .right({trees[93], lumberyards[93]}), .bottom_left({trees[141], lumberyards[141]}), .bottom({trees[142], lumberyards[142]}), .bottom_right({trees[143], lumberyards[143]}), .init(2'b10), .state({trees[92], lumberyards[92]}));
acre acre_1_43 (.clk(clk), .en(en), .top_left({trees[42], lumberyards[42]}), .top({trees[43], lumberyards[43]}), .top_right({trees[44], lumberyards[44]}), .left({trees[92], lumberyards[92]}), .right({trees[94], lumberyards[94]}), .bottom_left({trees[142], lumberyards[142]}), .bottom({trees[143], lumberyards[143]}), .bottom_right({trees[144], lumberyards[144]}), .init(2'b01), .state({trees[93], lumberyards[93]}));
acre acre_1_44 (.clk(clk), .en(en), .top_left({trees[43], lumberyards[43]}), .top({trees[44], lumberyards[44]}), .top_right({trees[45], lumberyards[45]}), .left({trees[93], lumberyards[93]}), .right({trees[95], lumberyards[95]}), .bottom_left({trees[143], lumberyards[143]}), .bottom({trees[144], lumberyards[144]}), .bottom_right({trees[145], lumberyards[145]}), .init(2'b10), .state({trees[94], lumberyards[94]}));
acre acre_1_45 (.clk(clk), .en(en), .top_left({trees[44], lumberyards[44]}), .top({trees[45], lumberyards[45]}), .top_right({trees[46], lumberyards[46]}), .left({trees[94], lumberyards[94]}), .right({trees[96], lumberyards[96]}), .bottom_left({trees[144], lumberyards[144]}), .bottom({trees[145], lumberyards[145]}), .bottom_right({trees[146], lumberyards[146]}), .init(2'b00), .state({trees[95], lumberyards[95]}));
acre acre_1_46 (.clk(clk), .en(en), .top_left({trees[45], lumberyards[45]}), .top({trees[46], lumberyards[46]}), .top_right({trees[47], lumberyards[47]}), .left({trees[95], lumberyards[95]}), .right({trees[97], lumberyards[97]}), .bottom_left({trees[145], lumberyards[145]}), .bottom({trees[146], lumberyards[146]}), .bottom_right({trees[147], lumberyards[147]}), .init(2'b00), .state({trees[96], lumberyards[96]}));
acre acre_1_47 (.clk(clk), .en(en), .top_left({trees[46], lumberyards[46]}), .top({trees[47], lumberyards[47]}), .top_right({trees[48], lumberyards[48]}), .left({trees[96], lumberyards[96]}), .right({trees[98], lumberyards[98]}), .bottom_left({trees[146], lumberyards[146]}), .bottom({trees[147], lumberyards[147]}), .bottom_right({trees[148], lumberyards[148]}), .init(2'b10), .state({trees[97], lumberyards[97]}));
acre acre_1_48 (.clk(clk), .en(en), .top_left({trees[47], lumberyards[47]}), .top({trees[48], lumberyards[48]}), .top_right({trees[49], lumberyards[49]}), .left({trees[97], lumberyards[97]}), .right({trees[99], lumberyards[99]}), .bottom_left({trees[147], lumberyards[147]}), .bottom({trees[148], lumberyards[148]}), .bottom_right({trees[149], lumberyards[149]}), .init(2'b00), .state({trees[98], lumberyards[98]}));
acre acre_1_49 (.clk(clk), .en(en), .top_left({trees[48], lumberyards[48]}), .top({trees[49], lumberyards[49]}), .top_right(2'b0), .left({trees[98], lumberyards[98]}), .right(2'b0), .bottom_left({trees[148], lumberyards[148]}), .bottom({trees[149], lumberyards[149]}), .bottom_right(2'b0), .init(2'b00), .state({trees[99], lumberyards[99]}));
acre acre_2_0 (.clk(clk), .en(en), .top_left(2'b0), .top({trees[50], lumberyards[50]}), .top_right({trees[51], lumberyards[51]}), .left(2'b0), .right({trees[101], lumberyards[101]}), .bottom_left(2'b0), .bottom({trees[150], lumberyards[150]}), .bottom_right({trees[151], lumberyards[151]}), .init(2'b01), .state({trees[100], lumberyards[100]}));
acre acre_2_1 (.clk(clk), .en(en), .top_left({trees[50], lumberyards[50]}), .top({trees[51], lumberyards[51]}), .top_right({trees[52], lumberyards[52]}), .left({trees[100], lumberyards[100]}), .right({trees[102], lumberyards[102]}), .bottom_left({trees[150], lumberyards[150]}), .bottom({trees[151], lumberyards[151]}), .bottom_right({trees[152], lumberyards[152]}), .init(2'b10), .state({trees[101], lumberyards[101]}));
acre acre_2_2 (.clk(clk), .en(en), .top_left({trees[51], lumberyards[51]}), .top({trees[52], lumberyards[52]}), .top_right({trees[53], lumberyards[53]}), .left({trees[101], lumberyards[101]}), .right({trees[103], lumberyards[103]}), .bottom_left({trees[151], lumberyards[151]}), .bottom({trees[152], lumberyards[152]}), .bottom_right({trees[153], lumberyards[153]}), .init(2'b00), .state({trees[102], lumberyards[102]}));
acre acre_2_3 (.clk(clk), .en(en), .top_left({trees[52], lumberyards[52]}), .top({trees[53], lumberyards[53]}), .top_right({trees[54], lumberyards[54]}), .left({trees[102], lumberyards[102]}), .right({trees[104], lumberyards[104]}), .bottom_left({trees[152], lumberyards[152]}), .bottom({trees[153], lumberyards[153]}), .bottom_right({trees[154], lumberyards[154]}), .init(2'b00), .state({trees[103], lumberyards[103]}));
acre acre_2_4 (.clk(clk), .en(en), .top_left({trees[53], lumberyards[53]}), .top({trees[54], lumberyards[54]}), .top_right({trees[55], lumberyards[55]}), .left({trees[103], lumberyards[103]}), .right({trees[105], lumberyards[105]}), .bottom_left({trees[153], lumberyards[153]}), .bottom({trees[154], lumberyards[154]}), .bottom_right({trees[155], lumberyards[155]}), .init(2'b00), .state({trees[104], lumberyards[104]}));
acre acre_2_5 (.clk(clk), .en(en), .top_left({trees[54], lumberyards[54]}), .top({trees[55], lumberyards[55]}), .top_right({trees[56], lumberyards[56]}), .left({trees[104], lumberyards[104]}), .right({trees[106], lumberyards[106]}), .bottom_left({trees[154], lumberyards[154]}), .bottom({trees[155], lumberyards[155]}), .bottom_right({trees[156], lumberyards[156]}), .init(2'b10), .state({trees[105], lumberyards[105]}));
acre acre_2_6 (.clk(clk), .en(en), .top_left({trees[55], lumberyards[55]}), .top({trees[56], lumberyards[56]}), .top_right({trees[57], lumberyards[57]}), .left({trees[105], lumberyards[105]}), .right({trees[107], lumberyards[107]}), .bottom_left({trees[155], lumberyards[155]}), .bottom({trees[156], lumberyards[156]}), .bottom_right({trees[157], lumberyards[157]}), .init(2'b00), .state({trees[106], lumberyards[106]}));
acre acre_2_7 (.clk(clk), .en(en), .top_left({trees[56], lumberyards[56]}), .top({trees[57], lumberyards[57]}), .top_right({trees[58], lumberyards[58]}), .left({trees[106], lumberyards[106]}), .right({trees[108], lumberyards[108]}), .bottom_left({trees[156], lumberyards[156]}), .bottom({trees[157], lumberyards[157]}), .bottom_right({trees[158], lumberyards[158]}), .init(2'b10), .state({trees[107], lumberyards[107]}));
acre acre_2_8 (.clk(clk), .en(en), .top_left({trees[57], lumberyards[57]}), .top({trees[58], lumberyards[58]}), .top_right({trees[59], lumberyards[59]}), .left({trees[107], lumberyards[107]}), .right({trees[109], lumberyards[109]}), .bottom_left({trees[157], lumberyards[157]}), .bottom({trees[158], lumberyards[158]}), .bottom_right({trees[159], lumberyards[159]}), .init(2'b00), .state({trees[108], lumberyards[108]}));
acre acre_2_9 (.clk(clk), .en(en), .top_left({trees[58], lumberyards[58]}), .top({trees[59], lumberyards[59]}), .top_right({trees[60], lumberyards[60]}), .left({trees[108], lumberyards[108]}), .right({trees[110], lumberyards[110]}), .bottom_left({trees[158], lumberyards[158]}), .bottom({trees[159], lumberyards[159]}), .bottom_right({trees[160], lumberyards[160]}), .init(2'b01), .state({trees[109], lumberyards[109]}));
acre acre_2_10 (.clk(clk), .en(en), .top_left({trees[59], lumberyards[59]}), .top({trees[60], lumberyards[60]}), .top_right({trees[61], lumberyards[61]}), .left({trees[109], lumberyards[109]}), .right({trees[111], lumberyards[111]}), .bottom_left({trees[159], lumberyards[159]}), .bottom({trees[160], lumberyards[160]}), .bottom_right({trees[161], lumberyards[161]}), .init(2'b00), .state({trees[110], lumberyards[110]}));
acre acre_2_11 (.clk(clk), .en(en), .top_left({trees[60], lumberyards[60]}), .top({trees[61], lumberyards[61]}), .top_right({trees[62], lumberyards[62]}), .left({trees[110], lumberyards[110]}), .right({trees[112], lumberyards[112]}), .bottom_left({trees[160], lumberyards[160]}), .bottom({trees[161], lumberyards[161]}), .bottom_right({trees[162], lumberyards[162]}), .init(2'b00), .state({trees[111], lumberyards[111]}));
acre acre_2_12 (.clk(clk), .en(en), .top_left({trees[61], lumberyards[61]}), .top({trees[62], lumberyards[62]}), .top_right({trees[63], lumberyards[63]}), .left({trees[111], lumberyards[111]}), .right({trees[113], lumberyards[113]}), .bottom_left({trees[161], lumberyards[161]}), .bottom({trees[162], lumberyards[162]}), .bottom_right({trees[163], lumberyards[163]}), .init(2'b10), .state({trees[112], lumberyards[112]}));
acre acre_2_13 (.clk(clk), .en(en), .top_left({trees[62], lumberyards[62]}), .top({trees[63], lumberyards[63]}), .top_right({trees[64], lumberyards[64]}), .left({trees[112], lumberyards[112]}), .right({trees[114], lumberyards[114]}), .bottom_left({trees[162], lumberyards[162]}), .bottom({trees[163], lumberyards[163]}), .bottom_right({trees[164], lumberyards[164]}), .init(2'b10), .state({trees[113], lumberyards[113]}));
acre acre_2_14 (.clk(clk), .en(en), .top_left({trees[63], lumberyards[63]}), .top({trees[64], lumberyards[64]}), .top_right({trees[65], lumberyards[65]}), .left({trees[113], lumberyards[113]}), .right({trees[115], lumberyards[115]}), .bottom_left({trees[163], lumberyards[163]}), .bottom({trees[164], lumberyards[164]}), .bottom_right({trees[165], lumberyards[165]}), .init(2'b00), .state({trees[114], lumberyards[114]}));
acre acre_2_15 (.clk(clk), .en(en), .top_left({trees[64], lumberyards[64]}), .top({trees[65], lumberyards[65]}), .top_right({trees[66], lumberyards[66]}), .left({trees[114], lumberyards[114]}), .right({trees[116], lumberyards[116]}), .bottom_left({trees[164], lumberyards[164]}), .bottom({trees[165], lumberyards[165]}), .bottom_right({trees[166], lumberyards[166]}), .init(2'b00), .state({trees[115], lumberyards[115]}));
acre acre_2_16 (.clk(clk), .en(en), .top_left({trees[65], lumberyards[65]}), .top({trees[66], lumberyards[66]}), .top_right({trees[67], lumberyards[67]}), .left({trees[115], lumberyards[115]}), .right({trees[117], lumberyards[117]}), .bottom_left({trees[165], lumberyards[165]}), .bottom({trees[166], lumberyards[166]}), .bottom_right({trees[167], lumberyards[167]}), .init(2'b00), .state({trees[116], lumberyards[116]}));
acre acre_2_17 (.clk(clk), .en(en), .top_left({trees[66], lumberyards[66]}), .top({trees[67], lumberyards[67]}), .top_right({trees[68], lumberyards[68]}), .left({trees[116], lumberyards[116]}), .right({trees[118], lumberyards[118]}), .bottom_left({trees[166], lumberyards[166]}), .bottom({trees[167], lumberyards[167]}), .bottom_right({trees[168], lumberyards[168]}), .init(2'b01), .state({trees[117], lumberyards[117]}));
acre acre_2_18 (.clk(clk), .en(en), .top_left({trees[67], lumberyards[67]}), .top({trees[68], lumberyards[68]}), .top_right({trees[69], lumberyards[69]}), .left({trees[117], lumberyards[117]}), .right({trees[119], lumberyards[119]}), .bottom_left({trees[167], lumberyards[167]}), .bottom({trees[168], lumberyards[168]}), .bottom_right({trees[169], lumberyards[169]}), .init(2'b10), .state({trees[118], lumberyards[118]}));
acre acre_2_19 (.clk(clk), .en(en), .top_left({trees[68], lumberyards[68]}), .top({trees[69], lumberyards[69]}), .top_right({trees[70], lumberyards[70]}), .left({trees[118], lumberyards[118]}), .right({trees[120], lumberyards[120]}), .bottom_left({trees[168], lumberyards[168]}), .bottom({trees[169], lumberyards[169]}), .bottom_right({trees[170], lumberyards[170]}), .init(2'b10), .state({trees[119], lumberyards[119]}));
acre acre_2_20 (.clk(clk), .en(en), .top_left({trees[69], lumberyards[69]}), .top({trees[70], lumberyards[70]}), .top_right({trees[71], lumberyards[71]}), .left({trees[119], lumberyards[119]}), .right({trees[121], lumberyards[121]}), .bottom_left({trees[169], lumberyards[169]}), .bottom({trees[170], lumberyards[170]}), .bottom_right({trees[171], lumberyards[171]}), .init(2'b10), .state({trees[120], lumberyards[120]}));
acre acre_2_21 (.clk(clk), .en(en), .top_left({trees[70], lumberyards[70]}), .top({trees[71], lumberyards[71]}), .top_right({trees[72], lumberyards[72]}), .left({trees[120], lumberyards[120]}), .right({trees[122], lumberyards[122]}), .bottom_left({trees[170], lumberyards[170]}), .bottom({trees[171], lumberyards[171]}), .bottom_right({trees[172], lumberyards[172]}), .init(2'b00), .state({trees[121], lumberyards[121]}));
acre acre_2_22 (.clk(clk), .en(en), .top_left({trees[71], lumberyards[71]}), .top({trees[72], lumberyards[72]}), .top_right({trees[73], lumberyards[73]}), .left({trees[121], lumberyards[121]}), .right({trees[123], lumberyards[123]}), .bottom_left({trees[171], lumberyards[171]}), .bottom({trees[172], lumberyards[172]}), .bottom_right({trees[173], lumberyards[173]}), .init(2'b00), .state({trees[122], lumberyards[122]}));
acre acre_2_23 (.clk(clk), .en(en), .top_left({trees[72], lumberyards[72]}), .top({trees[73], lumberyards[73]}), .top_right({trees[74], lumberyards[74]}), .left({trees[122], lumberyards[122]}), .right({trees[124], lumberyards[124]}), .bottom_left({trees[172], lumberyards[172]}), .bottom({trees[173], lumberyards[173]}), .bottom_right({trees[174], lumberyards[174]}), .init(2'b01), .state({trees[123], lumberyards[123]}));
acre acre_2_24 (.clk(clk), .en(en), .top_left({trees[73], lumberyards[73]}), .top({trees[74], lumberyards[74]}), .top_right({trees[75], lumberyards[75]}), .left({trees[123], lumberyards[123]}), .right({trees[125], lumberyards[125]}), .bottom_left({trees[173], lumberyards[173]}), .bottom({trees[174], lumberyards[174]}), .bottom_right({trees[175], lumberyards[175]}), .init(2'b10), .state({trees[124], lumberyards[124]}));
acre acre_2_25 (.clk(clk), .en(en), .top_left({trees[74], lumberyards[74]}), .top({trees[75], lumberyards[75]}), .top_right({trees[76], lumberyards[76]}), .left({trees[124], lumberyards[124]}), .right({trees[126], lumberyards[126]}), .bottom_left({trees[174], lumberyards[174]}), .bottom({trees[175], lumberyards[175]}), .bottom_right({trees[176], lumberyards[176]}), .init(2'b01), .state({trees[125], lumberyards[125]}));
acre acre_2_26 (.clk(clk), .en(en), .top_left({trees[75], lumberyards[75]}), .top({trees[76], lumberyards[76]}), .top_right({trees[77], lumberyards[77]}), .left({trees[125], lumberyards[125]}), .right({trees[127], lumberyards[127]}), .bottom_left({trees[175], lumberyards[175]}), .bottom({trees[176], lumberyards[176]}), .bottom_right({trees[177], lumberyards[177]}), .init(2'b00), .state({trees[126], lumberyards[126]}));
acre acre_2_27 (.clk(clk), .en(en), .top_left({trees[76], lumberyards[76]}), .top({trees[77], lumberyards[77]}), .top_right({trees[78], lumberyards[78]}), .left({trees[126], lumberyards[126]}), .right({trees[128], lumberyards[128]}), .bottom_left({trees[176], lumberyards[176]}), .bottom({trees[177], lumberyards[177]}), .bottom_right({trees[178], lumberyards[178]}), .init(2'b00), .state({trees[127], lumberyards[127]}));
acre acre_2_28 (.clk(clk), .en(en), .top_left({trees[77], lumberyards[77]}), .top({trees[78], lumberyards[78]}), .top_right({trees[79], lumberyards[79]}), .left({trees[127], lumberyards[127]}), .right({trees[129], lumberyards[129]}), .bottom_left({trees[177], lumberyards[177]}), .bottom({trees[178], lumberyards[178]}), .bottom_right({trees[179], lumberyards[179]}), .init(2'b01), .state({trees[128], lumberyards[128]}));
acre acre_2_29 (.clk(clk), .en(en), .top_left({trees[78], lumberyards[78]}), .top({trees[79], lumberyards[79]}), .top_right({trees[80], lumberyards[80]}), .left({trees[128], lumberyards[128]}), .right({trees[130], lumberyards[130]}), .bottom_left({trees[178], lumberyards[178]}), .bottom({trees[179], lumberyards[179]}), .bottom_right({trees[180], lumberyards[180]}), .init(2'b00), .state({trees[129], lumberyards[129]}));
acre acre_2_30 (.clk(clk), .en(en), .top_left({trees[79], lumberyards[79]}), .top({trees[80], lumberyards[80]}), .top_right({trees[81], lumberyards[81]}), .left({trees[129], lumberyards[129]}), .right({trees[131], lumberyards[131]}), .bottom_left({trees[179], lumberyards[179]}), .bottom({trees[180], lumberyards[180]}), .bottom_right({trees[181], lumberyards[181]}), .init(2'b00), .state({trees[130], lumberyards[130]}));
acre acre_2_31 (.clk(clk), .en(en), .top_left({trees[80], lumberyards[80]}), .top({trees[81], lumberyards[81]}), .top_right({trees[82], lumberyards[82]}), .left({trees[130], lumberyards[130]}), .right({trees[132], lumberyards[132]}), .bottom_left({trees[180], lumberyards[180]}), .bottom({trees[181], lumberyards[181]}), .bottom_right({trees[182], lumberyards[182]}), .init(2'b10), .state({trees[131], lumberyards[131]}));
acre acre_2_32 (.clk(clk), .en(en), .top_left({trees[81], lumberyards[81]}), .top({trees[82], lumberyards[82]}), .top_right({trees[83], lumberyards[83]}), .left({trees[131], lumberyards[131]}), .right({trees[133], lumberyards[133]}), .bottom_left({trees[181], lumberyards[181]}), .bottom({trees[182], lumberyards[182]}), .bottom_right({trees[183], lumberyards[183]}), .init(2'b00), .state({trees[132], lumberyards[132]}));
acre acre_2_33 (.clk(clk), .en(en), .top_left({trees[82], lumberyards[82]}), .top({trees[83], lumberyards[83]}), .top_right({trees[84], lumberyards[84]}), .left({trees[132], lumberyards[132]}), .right({trees[134], lumberyards[134]}), .bottom_left({trees[182], lumberyards[182]}), .bottom({trees[183], lumberyards[183]}), .bottom_right({trees[184], lumberyards[184]}), .init(2'b00), .state({trees[133], lumberyards[133]}));
acre acre_2_34 (.clk(clk), .en(en), .top_left({trees[83], lumberyards[83]}), .top({trees[84], lumberyards[84]}), .top_right({trees[85], lumberyards[85]}), .left({trees[133], lumberyards[133]}), .right({trees[135], lumberyards[135]}), .bottom_left({trees[183], lumberyards[183]}), .bottom({trees[184], lumberyards[184]}), .bottom_right({trees[185], lumberyards[185]}), .init(2'b00), .state({trees[134], lumberyards[134]}));
acre acre_2_35 (.clk(clk), .en(en), .top_left({trees[84], lumberyards[84]}), .top({trees[85], lumberyards[85]}), .top_right({trees[86], lumberyards[86]}), .left({trees[134], lumberyards[134]}), .right({trees[136], lumberyards[136]}), .bottom_left({trees[184], lumberyards[184]}), .bottom({trees[185], lumberyards[185]}), .bottom_right({trees[186], lumberyards[186]}), .init(2'b01), .state({trees[135], lumberyards[135]}));
acre acre_2_36 (.clk(clk), .en(en), .top_left({trees[85], lumberyards[85]}), .top({trees[86], lumberyards[86]}), .top_right({trees[87], lumberyards[87]}), .left({trees[135], lumberyards[135]}), .right({trees[137], lumberyards[137]}), .bottom_left({trees[185], lumberyards[185]}), .bottom({trees[186], lumberyards[186]}), .bottom_right({trees[187], lumberyards[187]}), .init(2'b00), .state({trees[136], lumberyards[136]}));
acre acre_2_37 (.clk(clk), .en(en), .top_left({trees[86], lumberyards[86]}), .top({trees[87], lumberyards[87]}), .top_right({trees[88], lumberyards[88]}), .left({trees[136], lumberyards[136]}), .right({trees[138], lumberyards[138]}), .bottom_left({trees[186], lumberyards[186]}), .bottom({trees[187], lumberyards[187]}), .bottom_right({trees[188], lumberyards[188]}), .init(2'b01), .state({trees[137], lumberyards[137]}));
acre acre_2_38 (.clk(clk), .en(en), .top_left({trees[87], lumberyards[87]}), .top({trees[88], lumberyards[88]}), .top_right({trees[89], lumberyards[89]}), .left({trees[137], lumberyards[137]}), .right({trees[139], lumberyards[139]}), .bottom_left({trees[187], lumberyards[187]}), .bottom({trees[188], lumberyards[188]}), .bottom_right({trees[189], lumberyards[189]}), .init(2'b01), .state({trees[138], lumberyards[138]}));
acre acre_2_39 (.clk(clk), .en(en), .top_left({trees[88], lumberyards[88]}), .top({trees[89], lumberyards[89]}), .top_right({trees[90], lumberyards[90]}), .left({trees[138], lumberyards[138]}), .right({trees[140], lumberyards[140]}), .bottom_left({trees[188], lumberyards[188]}), .bottom({trees[189], lumberyards[189]}), .bottom_right({trees[190], lumberyards[190]}), .init(2'b00), .state({trees[139], lumberyards[139]}));
acre acre_2_40 (.clk(clk), .en(en), .top_left({trees[89], lumberyards[89]}), .top({trees[90], lumberyards[90]}), .top_right({trees[91], lumberyards[91]}), .left({trees[139], lumberyards[139]}), .right({trees[141], lumberyards[141]}), .bottom_left({trees[189], lumberyards[189]}), .bottom({trees[190], lumberyards[190]}), .bottom_right({trees[191], lumberyards[191]}), .init(2'b10), .state({trees[140], lumberyards[140]}));
acre acre_2_41 (.clk(clk), .en(en), .top_left({trees[90], lumberyards[90]}), .top({trees[91], lumberyards[91]}), .top_right({trees[92], lumberyards[92]}), .left({trees[140], lumberyards[140]}), .right({trees[142], lumberyards[142]}), .bottom_left({trees[190], lumberyards[190]}), .bottom({trees[191], lumberyards[191]}), .bottom_right({trees[192], lumberyards[192]}), .init(2'b01), .state({trees[141], lumberyards[141]}));
acre acre_2_42 (.clk(clk), .en(en), .top_left({trees[91], lumberyards[91]}), .top({trees[92], lumberyards[92]}), .top_right({trees[93], lumberyards[93]}), .left({trees[141], lumberyards[141]}), .right({trees[143], lumberyards[143]}), .bottom_left({trees[191], lumberyards[191]}), .bottom({trees[192], lumberyards[192]}), .bottom_right({trees[193], lumberyards[193]}), .init(2'b01), .state({trees[142], lumberyards[142]}));
acre acre_2_43 (.clk(clk), .en(en), .top_left({trees[92], lumberyards[92]}), .top({trees[93], lumberyards[93]}), .top_right({trees[94], lumberyards[94]}), .left({trees[142], lumberyards[142]}), .right({trees[144], lumberyards[144]}), .bottom_left({trees[192], lumberyards[192]}), .bottom({trees[193], lumberyards[193]}), .bottom_right({trees[194], lumberyards[194]}), .init(2'b00), .state({trees[143], lumberyards[143]}));
acre acre_2_44 (.clk(clk), .en(en), .top_left({trees[93], lumberyards[93]}), .top({trees[94], lumberyards[94]}), .top_right({trees[95], lumberyards[95]}), .left({trees[143], lumberyards[143]}), .right({trees[145], lumberyards[145]}), .bottom_left({trees[193], lumberyards[193]}), .bottom({trees[194], lumberyards[194]}), .bottom_right({trees[195], lumberyards[195]}), .init(2'b00), .state({trees[144], lumberyards[144]}));
acre acre_2_45 (.clk(clk), .en(en), .top_left({trees[94], lumberyards[94]}), .top({trees[95], lumberyards[95]}), .top_right({trees[96], lumberyards[96]}), .left({trees[144], lumberyards[144]}), .right({trees[146], lumberyards[146]}), .bottom_left({trees[194], lumberyards[194]}), .bottom({trees[195], lumberyards[195]}), .bottom_right({trees[196], lumberyards[196]}), .init(2'b00), .state({trees[145], lumberyards[145]}));
acre acre_2_46 (.clk(clk), .en(en), .top_left({trees[95], lumberyards[95]}), .top({trees[96], lumberyards[96]}), .top_right({trees[97], lumberyards[97]}), .left({trees[145], lumberyards[145]}), .right({trees[147], lumberyards[147]}), .bottom_left({trees[195], lumberyards[195]}), .bottom({trees[196], lumberyards[196]}), .bottom_right({trees[197], lumberyards[197]}), .init(2'b00), .state({trees[146], lumberyards[146]}));
acre acre_2_47 (.clk(clk), .en(en), .top_left({trees[96], lumberyards[96]}), .top({trees[97], lumberyards[97]}), .top_right({trees[98], lumberyards[98]}), .left({trees[146], lumberyards[146]}), .right({trees[148], lumberyards[148]}), .bottom_left({trees[196], lumberyards[196]}), .bottom({trees[197], lumberyards[197]}), .bottom_right({trees[198], lumberyards[198]}), .init(2'b00), .state({trees[147], lumberyards[147]}));
acre acre_2_48 (.clk(clk), .en(en), .top_left({trees[97], lumberyards[97]}), .top({trees[98], lumberyards[98]}), .top_right({trees[99], lumberyards[99]}), .left({trees[147], lumberyards[147]}), .right({trees[149], lumberyards[149]}), .bottom_left({trees[197], lumberyards[197]}), .bottom({trees[198], lumberyards[198]}), .bottom_right({trees[199], lumberyards[199]}), .init(2'b00), .state({trees[148], lumberyards[148]}));
acre acre_2_49 (.clk(clk), .en(en), .top_left({trees[98], lumberyards[98]}), .top({trees[99], lumberyards[99]}), .top_right(2'b0), .left({trees[148], lumberyards[148]}), .right(2'b0), .bottom_left({trees[198], lumberyards[198]}), .bottom({trees[199], lumberyards[199]}), .bottom_right(2'b0), .init(2'b00), .state({trees[149], lumberyards[149]}));
acre acre_3_0 (.clk(clk), .en(en), .top_left(2'b0), .top({trees[100], lumberyards[100]}), .top_right({trees[101], lumberyards[101]}), .left(2'b0), .right({trees[151], lumberyards[151]}), .bottom_left(2'b0), .bottom({trees[200], lumberyards[200]}), .bottom_right({trees[201], lumberyards[201]}), .init(2'b01), .state({trees[150], lumberyards[150]}));
acre acre_3_1 (.clk(clk), .en(en), .top_left({trees[100], lumberyards[100]}), .top({trees[101], lumberyards[101]}), .top_right({trees[102], lumberyards[102]}), .left({trees[150], lumberyards[150]}), .right({trees[152], lumberyards[152]}), .bottom_left({trees[200], lumberyards[200]}), .bottom({trees[201], lumberyards[201]}), .bottom_right({trees[202], lumberyards[202]}), .init(2'b01), .state({trees[151], lumberyards[151]}));
acre acre_3_2 (.clk(clk), .en(en), .top_left({trees[101], lumberyards[101]}), .top({trees[102], lumberyards[102]}), .top_right({trees[103], lumberyards[103]}), .left({trees[151], lumberyards[151]}), .right({trees[153], lumberyards[153]}), .bottom_left({trees[201], lumberyards[201]}), .bottom({trees[202], lumberyards[202]}), .bottom_right({trees[203], lumberyards[203]}), .init(2'b00), .state({trees[152], lumberyards[152]}));
acre acre_3_3 (.clk(clk), .en(en), .top_left({trees[102], lumberyards[102]}), .top({trees[103], lumberyards[103]}), .top_right({trees[104], lumberyards[104]}), .left({trees[152], lumberyards[152]}), .right({trees[154], lumberyards[154]}), .bottom_left({trees[202], lumberyards[202]}), .bottom({trees[203], lumberyards[203]}), .bottom_right({trees[204], lumberyards[204]}), .init(2'b00), .state({trees[153], lumberyards[153]}));
acre acre_3_4 (.clk(clk), .en(en), .top_left({trees[103], lumberyards[103]}), .top({trees[104], lumberyards[104]}), .top_right({trees[105], lumberyards[105]}), .left({trees[153], lumberyards[153]}), .right({trees[155], lumberyards[155]}), .bottom_left({trees[203], lumberyards[203]}), .bottom({trees[204], lumberyards[204]}), .bottom_right({trees[205], lumberyards[205]}), .init(2'b00), .state({trees[154], lumberyards[154]}));
acre acre_3_5 (.clk(clk), .en(en), .top_left({trees[104], lumberyards[104]}), .top({trees[105], lumberyards[105]}), .top_right({trees[106], lumberyards[106]}), .left({trees[154], lumberyards[154]}), .right({trees[156], lumberyards[156]}), .bottom_left({trees[204], lumberyards[204]}), .bottom({trees[205], lumberyards[205]}), .bottom_right({trees[206], lumberyards[206]}), .init(2'b00), .state({trees[155], lumberyards[155]}));
acre acre_3_6 (.clk(clk), .en(en), .top_left({trees[105], lumberyards[105]}), .top({trees[106], lumberyards[106]}), .top_right({trees[107], lumberyards[107]}), .left({trees[155], lumberyards[155]}), .right({trees[157], lumberyards[157]}), .bottom_left({trees[205], lumberyards[205]}), .bottom({trees[206], lumberyards[206]}), .bottom_right({trees[207], lumberyards[207]}), .init(2'b00), .state({trees[156], lumberyards[156]}));
acre acre_3_7 (.clk(clk), .en(en), .top_left({trees[106], lumberyards[106]}), .top({trees[107], lumberyards[107]}), .top_right({trees[108], lumberyards[108]}), .left({trees[156], lumberyards[156]}), .right({trees[158], lumberyards[158]}), .bottom_left({trees[206], lumberyards[206]}), .bottom({trees[207], lumberyards[207]}), .bottom_right({trees[208], lumberyards[208]}), .init(2'b01), .state({trees[157], lumberyards[157]}));
acre acre_3_8 (.clk(clk), .en(en), .top_left({trees[107], lumberyards[107]}), .top({trees[108], lumberyards[108]}), .top_right({trees[109], lumberyards[109]}), .left({trees[157], lumberyards[157]}), .right({trees[159], lumberyards[159]}), .bottom_left({trees[207], lumberyards[207]}), .bottom({trees[208], lumberyards[208]}), .bottom_right({trees[209], lumberyards[209]}), .init(2'b00), .state({trees[158], lumberyards[158]}));
acre acre_3_9 (.clk(clk), .en(en), .top_left({trees[108], lumberyards[108]}), .top({trees[109], lumberyards[109]}), .top_right({trees[110], lumberyards[110]}), .left({trees[158], lumberyards[158]}), .right({trees[160], lumberyards[160]}), .bottom_left({trees[208], lumberyards[208]}), .bottom({trees[209], lumberyards[209]}), .bottom_right({trees[210], lumberyards[210]}), .init(2'b00), .state({trees[159], lumberyards[159]}));
acre acre_3_10 (.clk(clk), .en(en), .top_left({trees[109], lumberyards[109]}), .top({trees[110], lumberyards[110]}), .top_right({trees[111], lumberyards[111]}), .left({trees[159], lumberyards[159]}), .right({trees[161], lumberyards[161]}), .bottom_left({trees[209], lumberyards[209]}), .bottom({trees[210], lumberyards[210]}), .bottom_right({trees[211], lumberyards[211]}), .init(2'b10), .state({trees[160], lumberyards[160]}));
acre acre_3_11 (.clk(clk), .en(en), .top_left({trees[110], lumberyards[110]}), .top({trees[111], lumberyards[111]}), .top_right({trees[112], lumberyards[112]}), .left({trees[160], lumberyards[160]}), .right({trees[162], lumberyards[162]}), .bottom_left({trees[210], lumberyards[210]}), .bottom({trees[211], lumberyards[211]}), .bottom_right({trees[212], lumberyards[212]}), .init(2'b01), .state({trees[161], lumberyards[161]}));
acre acre_3_12 (.clk(clk), .en(en), .top_left({trees[111], lumberyards[111]}), .top({trees[112], lumberyards[112]}), .top_right({trees[113], lumberyards[113]}), .left({trees[161], lumberyards[161]}), .right({trees[163], lumberyards[163]}), .bottom_left({trees[211], lumberyards[211]}), .bottom({trees[212], lumberyards[212]}), .bottom_right({trees[213], lumberyards[213]}), .init(2'b00), .state({trees[162], lumberyards[162]}));
acre acre_3_13 (.clk(clk), .en(en), .top_left({trees[112], lumberyards[112]}), .top({trees[113], lumberyards[113]}), .top_right({trees[114], lumberyards[114]}), .left({trees[162], lumberyards[162]}), .right({trees[164], lumberyards[164]}), .bottom_left({trees[212], lumberyards[212]}), .bottom({trees[213], lumberyards[213]}), .bottom_right({trees[214], lumberyards[214]}), .init(2'b00), .state({trees[163], lumberyards[163]}));
acre acre_3_14 (.clk(clk), .en(en), .top_left({trees[113], lumberyards[113]}), .top({trees[114], lumberyards[114]}), .top_right({trees[115], lumberyards[115]}), .left({trees[163], lumberyards[163]}), .right({trees[165], lumberyards[165]}), .bottom_left({trees[213], lumberyards[213]}), .bottom({trees[214], lumberyards[214]}), .bottom_right({trees[215], lumberyards[215]}), .init(2'b00), .state({trees[164], lumberyards[164]}));
acre acre_3_15 (.clk(clk), .en(en), .top_left({trees[114], lumberyards[114]}), .top({trees[115], lumberyards[115]}), .top_right({trees[116], lumberyards[116]}), .left({trees[164], lumberyards[164]}), .right({trees[166], lumberyards[166]}), .bottom_left({trees[214], lumberyards[214]}), .bottom({trees[215], lumberyards[215]}), .bottom_right({trees[216], lumberyards[216]}), .init(2'b00), .state({trees[165], lumberyards[165]}));
acre acre_3_16 (.clk(clk), .en(en), .top_left({trees[115], lumberyards[115]}), .top({trees[116], lumberyards[116]}), .top_right({trees[117], lumberyards[117]}), .left({trees[165], lumberyards[165]}), .right({trees[167], lumberyards[167]}), .bottom_left({trees[215], lumberyards[215]}), .bottom({trees[216], lumberyards[216]}), .bottom_right({trees[217], lumberyards[217]}), .init(2'b00), .state({trees[166], lumberyards[166]}));
acre acre_3_17 (.clk(clk), .en(en), .top_left({trees[116], lumberyards[116]}), .top({trees[117], lumberyards[117]}), .top_right({trees[118], lumberyards[118]}), .left({trees[166], lumberyards[166]}), .right({trees[168], lumberyards[168]}), .bottom_left({trees[216], lumberyards[216]}), .bottom({trees[217], lumberyards[217]}), .bottom_right({trees[218], lumberyards[218]}), .init(2'b01), .state({trees[167], lumberyards[167]}));
acre acre_3_18 (.clk(clk), .en(en), .top_left({trees[117], lumberyards[117]}), .top({trees[118], lumberyards[118]}), .top_right({trees[119], lumberyards[119]}), .left({trees[167], lumberyards[167]}), .right({trees[169], lumberyards[169]}), .bottom_left({trees[217], lumberyards[217]}), .bottom({trees[218], lumberyards[218]}), .bottom_right({trees[219], lumberyards[219]}), .init(2'b00), .state({trees[168], lumberyards[168]}));
acre acre_3_19 (.clk(clk), .en(en), .top_left({trees[118], lumberyards[118]}), .top({trees[119], lumberyards[119]}), .top_right({trees[120], lumberyards[120]}), .left({trees[168], lumberyards[168]}), .right({trees[170], lumberyards[170]}), .bottom_left({trees[218], lumberyards[218]}), .bottom({trees[219], lumberyards[219]}), .bottom_right({trees[220], lumberyards[220]}), .init(2'b00), .state({trees[169], lumberyards[169]}));
acre acre_3_20 (.clk(clk), .en(en), .top_left({trees[119], lumberyards[119]}), .top({trees[120], lumberyards[120]}), .top_right({trees[121], lumberyards[121]}), .left({trees[169], lumberyards[169]}), .right({trees[171], lumberyards[171]}), .bottom_left({trees[219], lumberyards[219]}), .bottom({trees[220], lumberyards[220]}), .bottom_right({trees[221], lumberyards[221]}), .init(2'b00), .state({trees[170], lumberyards[170]}));
acre acre_3_21 (.clk(clk), .en(en), .top_left({trees[120], lumberyards[120]}), .top({trees[121], lumberyards[121]}), .top_right({trees[122], lumberyards[122]}), .left({trees[170], lumberyards[170]}), .right({trees[172], lumberyards[172]}), .bottom_left({trees[220], lumberyards[220]}), .bottom({trees[221], lumberyards[221]}), .bottom_right({trees[222], lumberyards[222]}), .init(2'b00), .state({trees[171], lumberyards[171]}));
acre acre_3_22 (.clk(clk), .en(en), .top_left({trees[121], lumberyards[121]}), .top({trees[122], lumberyards[122]}), .top_right({trees[123], lumberyards[123]}), .left({trees[171], lumberyards[171]}), .right({trees[173], lumberyards[173]}), .bottom_left({trees[221], lumberyards[221]}), .bottom({trees[222], lumberyards[222]}), .bottom_right({trees[223], lumberyards[223]}), .init(2'b00), .state({trees[172], lumberyards[172]}));
acre acre_3_23 (.clk(clk), .en(en), .top_left({trees[122], lumberyards[122]}), .top({trees[123], lumberyards[123]}), .top_right({trees[124], lumberyards[124]}), .left({trees[172], lumberyards[172]}), .right({trees[174], lumberyards[174]}), .bottom_left({trees[222], lumberyards[222]}), .bottom({trees[223], lumberyards[223]}), .bottom_right({trees[224], lumberyards[224]}), .init(2'b01), .state({trees[173], lumberyards[173]}));
acre acre_3_24 (.clk(clk), .en(en), .top_left({trees[123], lumberyards[123]}), .top({trees[124], lumberyards[124]}), .top_right({trees[125], lumberyards[125]}), .left({trees[173], lumberyards[173]}), .right({trees[175], lumberyards[175]}), .bottom_left({trees[223], lumberyards[223]}), .bottom({trees[224], lumberyards[224]}), .bottom_right({trees[225], lumberyards[225]}), .init(2'b00), .state({trees[174], lumberyards[174]}));
acre acre_3_25 (.clk(clk), .en(en), .top_left({trees[124], lumberyards[124]}), .top({trees[125], lumberyards[125]}), .top_right({trees[126], lumberyards[126]}), .left({trees[174], lumberyards[174]}), .right({trees[176], lumberyards[176]}), .bottom_left({trees[224], lumberyards[224]}), .bottom({trees[225], lumberyards[225]}), .bottom_right({trees[226], lumberyards[226]}), .init(2'b10), .state({trees[175], lumberyards[175]}));
acre acre_3_26 (.clk(clk), .en(en), .top_left({trees[125], lumberyards[125]}), .top({trees[126], lumberyards[126]}), .top_right({trees[127], lumberyards[127]}), .left({trees[175], lumberyards[175]}), .right({trees[177], lumberyards[177]}), .bottom_left({trees[225], lumberyards[225]}), .bottom({trees[226], lumberyards[226]}), .bottom_right({trees[227], lumberyards[227]}), .init(2'b00), .state({trees[176], lumberyards[176]}));
acre acre_3_27 (.clk(clk), .en(en), .top_left({trees[126], lumberyards[126]}), .top({trees[127], lumberyards[127]}), .top_right({trees[128], lumberyards[128]}), .left({trees[176], lumberyards[176]}), .right({trees[178], lumberyards[178]}), .bottom_left({trees[226], lumberyards[226]}), .bottom({trees[227], lumberyards[227]}), .bottom_right({trees[228], lumberyards[228]}), .init(2'b00), .state({trees[177], lumberyards[177]}));
acre acre_3_28 (.clk(clk), .en(en), .top_left({trees[127], lumberyards[127]}), .top({trees[128], lumberyards[128]}), .top_right({trees[129], lumberyards[129]}), .left({trees[177], lumberyards[177]}), .right({trees[179], lumberyards[179]}), .bottom_left({trees[227], lumberyards[227]}), .bottom({trees[228], lumberyards[228]}), .bottom_right({trees[229], lumberyards[229]}), .init(2'b00), .state({trees[178], lumberyards[178]}));
acre acre_3_29 (.clk(clk), .en(en), .top_left({trees[128], lumberyards[128]}), .top({trees[129], lumberyards[129]}), .top_right({trees[130], lumberyards[130]}), .left({trees[178], lumberyards[178]}), .right({trees[180], lumberyards[180]}), .bottom_left({trees[228], lumberyards[228]}), .bottom({trees[229], lumberyards[229]}), .bottom_right({trees[230], lumberyards[230]}), .init(2'b00), .state({trees[179], lumberyards[179]}));
acre acre_3_30 (.clk(clk), .en(en), .top_left({trees[129], lumberyards[129]}), .top({trees[130], lumberyards[130]}), .top_right({trees[131], lumberyards[131]}), .left({trees[179], lumberyards[179]}), .right({trees[181], lumberyards[181]}), .bottom_left({trees[229], lumberyards[229]}), .bottom({trees[230], lumberyards[230]}), .bottom_right({trees[231], lumberyards[231]}), .init(2'b01), .state({trees[180], lumberyards[180]}));
acre acre_3_31 (.clk(clk), .en(en), .top_left({trees[130], lumberyards[130]}), .top({trees[131], lumberyards[131]}), .top_right({trees[132], lumberyards[132]}), .left({trees[180], lumberyards[180]}), .right({trees[182], lumberyards[182]}), .bottom_left({trees[230], lumberyards[230]}), .bottom({trees[231], lumberyards[231]}), .bottom_right({trees[232], lumberyards[232]}), .init(2'b00), .state({trees[181], lumberyards[181]}));
acre acre_3_32 (.clk(clk), .en(en), .top_left({trees[131], lumberyards[131]}), .top({trees[132], lumberyards[132]}), .top_right({trees[133], lumberyards[133]}), .left({trees[181], lumberyards[181]}), .right({trees[183], lumberyards[183]}), .bottom_left({trees[231], lumberyards[231]}), .bottom({trees[232], lumberyards[232]}), .bottom_right({trees[233], lumberyards[233]}), .init(2'b00), .state({trees[182], lumberyards[182]}));
acre acre_3_33 (.clk(clk), .en(en), .top_left({trees[132], lumberyards[132]}), .top({trees[133], lumberyards[133]}), .top_right({trees[134], lumberyards[134]}), .left({trees[182], lumberyards[182]}), .right({trees[184], lumberyards[184]}), .bottom_left({trees[232], lumberyards[232]}), .bottom({trees[233], lumberyards[233]}), .bottom_right({trees[234], lumberyards[234]}), .init(2'b10), .state({trees[183], lumberyards[183]}));
acre acre_3_34 (.clk(clk), .en(en), .top_left({trees[133], lumberyards[133]}), .top({trees[134], lumberyards[134]}), .top_right({trees[135], lumberyards[135]}), .left({trees[183], lumberyards[183]}), .right({trees[185], lumberyards[185]}), .bottom_left({trees[233], lumberyards[233]}), .bottom({trees[234], lumberyards[234]}), .bottom_right({trees[235], lumberyards[235]}), .init(2'b00), .state({trees[184], lumberyards[184]}));
acre acre_3_35 (.clk(clk), .en(en), .top_left({trees[134], lumberyards[134]}), .top({trees[135], lumberyards[135]}), .top_right({trees[136], lumberyards[136]}), .left({trees[184], lumberyards[184]}), .right({trees[186], lumberyards[186]}), .bottom_left({trees[234], lumberyards[234]}), .bottom({trees[235], lumberyards[235]}), .bottom_right({trees[236], lumberyards[236]}), .init(2'b10), .state({trees[185], lumberyards[185]}));
acre acre_3_36 (.clk(clk), .en(en), .top_left({trees[135], lumberyards[135]}), .top({trees[136], lumberyards[136]}), .top_right({trees[137], lumberyards[137]}), .left({trees[185], lumberyards[185]}), .right({trees[187], lumberyards[187]}), .bottom_left({trees[235], lumberyards[235]}), .bottom({trees[236], lumberyards[236]}), .bottom_right({trees[237], lumberyards[237]}), .init(2'b01), .state({trees[186], lumberyards[186]}));
acre acre_3_37 (.clk(clk), .en(en), .top_left({trees[136], lumberyards[136]}), .top({trees[137], lumberyards[137]}), .top_right({trees[138], lumberyards[138]}), .left({trees[186], lumberyards[186]}), .right({trees[188], lumberyards[188]}), .bottom_left({trees[236], lumberyards[236]}), .bottom({trees[237], lumberyards[237]}), .bottom_right({trees[238], lumberyards[238]}), .init(2'b10), .state({trees[187], lumberyards[187]}));
acre acre_3_38 (.clk(clk), .en(en), .top_left({trees[137], lumberyards[137]}), .top({trees[138], lumberyards[138]}), .top_right({trees[139], lumberyards[139]}), .left({trees[187], lumberyards[187]}), .right({trees[189], lumberyards[189]}), .bottom_left({trees[237], lumberyards[237]}), .bottom({trees[238], lumberyards[238]}), .bottom_right({trees[239], lumberyards[239]}), .init(2'b00), .state({trees[188], lumberyards[188]}));
acre acre_3_39 (.clk(clk), .en(en), .top_left({trees[138], lumberyards[138]}), .top({trees[139], lumberyards[139]}), .top_right({trees[140], lumberyards[140]}), .left({trees[188], lumberyards[188]}), .right({trees[190], lumberyards[190]}), .bottom_left({trees[238], lumberyards[238]}), .bottom({trees[239], lumberyards[239]}), .bottom_right({trees[240], lumberyards[240]}), .init(2'b00), .state({trees[189], lumberyards[189]}));
acre acre_3_40 (.clk(clk), .en(en), .top_left({trees[139], lumberyards[139]}), .top({trees[140], lumberyards[140]}), .top_right({trees[141], lumberyards[141]}), .left({trees[189], lumberyards[189]}), .right({trees[191], lumberyards[191]}), .bottom_left({trees[239], lumberyards[239]}), .bottom({trees[240], lumberyards[240]}), .bottom_right({trees[241], lumberyards[241]}), .init(2'b00), .state({trees[190], lumberyards[190]}));
acre acre_3_41 (.clk(clk), .en(en), .top_left({trees[140], lumberyards[140]}), .top({trees[141], lumberyards[141]}), .top_right({trees[142], lumberyards[142]}), .left({trees[190], lumberyards[190]}), .right({trees[192], lumberyards[192]}), .bottom_left({trees[240], lumberyards[240]}), .bottom({trees[241], lumberyards[241]}), .bottom_right({trees[242], lumberyards[242]}), .init(2'b00), .state({trees[191], lumberyards[191]}));
acre acre_3_42 (.clk(clk), .en(en), .top_left({trees[141], lumberyards[141]}), .top({trees[142], lumberyards[142]}), .top_right({trees[143], lumberyards[143]}), .left({trees[191], lumberyards[191]}), .right({trees[193], lumberyards[193]}), .bottom_left({trees[241], lumberyards[241]}), .bottom({trees[242], lumberyards[242]}), .bottom_right({trees[243], lumberyards[243]}), .init(2'b10), .state({trees[192], lumberyards[192]}));
acre acre_3_43 (.clk(clk), .en(en), .top_left({trees[142], lumberyards[142]}), .top({trees[143], lumberyards[143]}), .top_right({trees[144], lumberyards[144]}), .left({trees[192], lumberyards[192]}), .right({trees[194], lumberyards[194]}), .bottom_left({trees[242], lumberyards[242]}), .bottom({trees[243], lumberyards[243]}), .bottom_right({trees[244], lumberyards[244]}), .init(2'b00), .state({trees[193], lumberyards[193]}));
acre acre_3_44 (.clk(clk), .en(en), .top_left({trees[143], lumberyards[143]}), .top({trees[144], lumberyards[144]}), .top_right({trees[145], lumberyards[145]}), .left({trees[193], lumberyards[193]}), .right({trees[195], lumberyards[195]}), .bottom_left({trees[243], lumberyards[243]}), .bottom({trees[244], lumberyards[244]}), .bottom_right({trees[245], lumberyards[245]}), .init(2'b00), .state({trees[194], lumberyards[194]}));
acre acre_3_45 (.clk(clk), .en(en), .top_left({trees[144], lumberyards[144]}), .top({trees[145], lumberyards[145]}), .top_right({trees[146], lumberyards[146]}), .left({trees[194], lumberyards[194]}), .right({trees[196], lumberyards[196]}), .bottom_left({trees[244], lumberyards[244]}), .bottom({trees[245], lumberyards[245]}), .bottom_right({trees[246], lumberyards[246]}), .init(2'b00), .state({trees[195], lumberyards[195]}));
acre acre_3_46 (.clk(clk), .en(en), .top_left({trees[145], lumberyards[145]}), .top({trees[146], lumberyards[146]}), .top_right({trees[147], lumberyards[147]}), .left({trees[195], lumberyards[195]}), .right({trees[197], lumberyards[197]}), .bottom_left({trees[245], lumberyards[245]}), .bottom({trees[246], lumberyards[246]}), .bottom_right({trees[247], lumberyards[247]}), .init(2'b01), .state({trees[196], lumberyards[196]}));
acre acre_3_47 (.clk(clk), .en(en), .top_left({trees[146], lumberyards[146]}), .top({trees[147], lumberyards[147]}), .top_right({trees[148], lumberyards[148]}), .left({trees[196], lumberyards[196]}), .right({trees[198], lumberyards[198]}), .bottom_left({trees[246], lumberyards[246]}), .bottom({trees[247], lumberyards[247]}), .bottom_right({trees[248], lumberyards[248]}), .init(2'b10), .state({trees[197], lumberyards[197]}));
acre acre_3_48 (.clk(clk), .en(en), .top_left({trees[147], lumberyards[147]}), .top({trees[148], lumberyards[148]}), .top_right({trees[149], lumberyards[149]}), .left({trees[197], lumberyards[197]}), .right({trees[199], lumberyards[199]}), .bottom_left({trees[247], lumberyards[247]}), .bottom({trees[248], lumberyards[248]}), .bottom_right({trees[249], lumberyards[249]}), .init(2'b00), .state({trees[198], lumberyards[198]}));
acre acre_3_49 (.clk(clk), .en(en), .top_left({trees[148], lumberyards[148]}), .top({trees[149], lumberyards[149]}), .top_right(2'b0), .left({trees[198], lumberyards[198]}), .right(2'b0), .bottom_left({trees[248], lumberyards[248]}), .bottom({trees[249], lumberyards[249]}), .bottom_right(2'b0), .init(2'b00), .state({trees[199], lumberyards[199]}));
acre acre_4_0 (.clk(clk), .en(en), .top_left(2'b0), .top({trees[150], lumberyards[150]}), .top_right({trees[151], lumberyards[151]}), .left(2'b0), .right({trees[201], lumberyards[201]}), .bottom_left(2'b0), .bottom({trees[250], lumberyards[250]}), .bottom_right({trees[251], lumberyards[251]}), .init(2'b01), .state({trees[200], lumberyards[200]}));
acre acre_4_1 (.clk(clk), .en(en), .top_left({trees[150], lumberyards[150]}), .top({trees[151], lumberyards[151]}), .top_right({trees[152], lumberyards[152]}), .left({trees[200], lumberyards[200]}), .right({trees[202], lumberyards[202]}), .bottom_left({trees[250], lumberyards[250]}), .bottom({trees[251], lumberyards[251]}), .bottom_right({trees[252], lumberyards[252]}), .init(2'b00), .state({trees[201], lumberyards[201]}));
acre acre_4_2 (.clk(clk), .en(en), .top_left({trees[151], lumberyards[151]}), .top({trees[152], lumberyards[152]}), .top_right({trees[153], lumberyards[153]}), .left({trees[201], lumberyards[201]}), .right({trees[203], lumberyards[203]}), .bottom_left({trees[251], lumberyards[251]}), .bottom({trees[252], lumberyards[252]}), .bottom_right({trees[253], lumberyards[253]}), .init(2'b00), .state({trees[202], lumberyards[202]}));
acre acre_4_3 (.clk(clk), .en(en), .top_left({trees[152], lumberyards[152]}), .top({trees[153], lumberyards[153]}), .top_right({trees[154], lumberyards[154]}), .left({trees[202], lumberyards[202]}), .right({trees[204], lumberyards[204]}), .bottom_left({trees[252], lumberyards[252]}), .bottom({trees[253], lumberyards[253]}), .bottom_right({trees[254], lumberyards[254]}), .init(2'b00), .state({trees[203], lumberyards[203]}));
acre acre_4_4 (.clk(clk), .en(en), .top_left({trees[153], lumberyards[153]}), .top({trees[154], lumberyards[154]}), .top_right({trees[155], lumberyards[155]}), .left({trees[203], lumberyards[203]}), .right({trees[205], lumberyards[205]}), .bottom_left({trees[253], lumberyards[253]}), .bottom({trees[254], lumberyards[254]}), .bottom_right({trees[255], lumberyards[255]}), .init(2'b00), .state({trees[204], lumberyards[204]}));
acre acre_4_5 (.clk(clk), .en(en), .top_left({trees[154], lumberyards[154]}), .top({trees[155], lumberyards[155]}), .top_right({trees[156], lumberyards[156]}), .left({trees[204], lumberyards[204]}), .right({trees[206], lumberyards[206]}), .bottom_left({trees[254], lumberyards[254]}), .bottom({trees[255], lumberyards[255]}), .bottom_right({trees[256], lumberyards[256]}), .init(2'b10), .state({trees[205], lumberyards[205]}));
acre acre_4_6 (.clk(clk), .en(en), .top_left({trees[155], lumberyards[155]}), .top({trees[156], lumberyards[156]}), .top_right({trees[157], lumberyards[157]}), .left({trees[205], lumberyards[205]}), .right({trees[207], lumberyards[207]}), .bottom_left({trees[255], lumberyards[255]}), .bottom({trees[256], lumberyards[256]}), .bottom_right({trees[257], lumberyards[257]}), .init(2'b00), .state({trees[206], lumberyards[206]}));
acre acre_4_7 (.clk(clk), .en(en), .top_left({trees[156], lumberyards[156]}), .top({trees[157], lumberyards[157]}), .top_right({trees[158], lumberyards[158]}), .left({trees[206], lumberyards[206]}), .right({trees[208], lumberyards[208]}), .bottom_left({trees[256], lumberyards[256]}), .bottom({trees[257], lumberyards[257]}), .bottom_right({trees[258], lumberyards[258]}), .init(2'b00), .state({trees[207], lumberyards[207]}));
acre acre_4_8 (.clk(clk), .en(en), .top_left({trees[157], lumberyards[157]}), .top({trees[158], lumberyards[158]}), .top_right({trees[159], lumberyards[159]}), .left({trees[207], lumberyards[207]}), .right({trees[209], lumberyards[209]}), .bottom_left({trees[257], lumberyards[257]}), .bottom({trees[258], lumberyards[258]}), .bottom_right({trees[259], lumberyards[259]}), .init(2'b00), .state({trees[208], lumberyards[208]}));
acre acre_4_9 (.clk(clk), .en(en), .top_left({trees[158], lumberyards[158]}), .top({trees[159], lumberyards[159]}), .top_right({trees[160], lumberyards[160]}), .left({trees[208], lumberyards[208]}), .right({trees[210], lumberyards[210]}), .bottom_left({trees[258], lumberyards[258]}), .bottom({trees[259], lumberyards[259]}), .bottom_right({trees[260], lumberyards[260]}), .init(2'b00), .state({trees[209], lumberyards[209]}));
acre acre_4_10 (.clk(clk), .en(en), .top_left({trees[159], lumberyards[159]}), .top({trees[160], lumberyards[160]}), .top_right({trees[161], lumberyards[161]}), .left({trees[209], lumberyards[209]}), .right({trees[211], lumberyards[211]}), .bottom_left({trees[259], lumberyards[259]}), .bottom({trees[260], lumberyards[260]}), .bottom_right({trees[261], lumberyards[261]}), .init(2'b00), .state({trees[210], lumberyards[210]}));
acre acre_4_11 (.clk(clk), .en(en), .top_left({trees[160], lumberyards[160]}), .top({trees[161], lumberyards[161]}), .top_right({trees[162], lumberyards[162]}), .left({trees[210], lumberyards[210]}), .right({trees[212], lumberyards[212]}), .bottom_left({trees[260], lumberyards[260]}), .bottom({trees[261], lumberyards[261]}), .bottom_right({trees[262], lumberyards[262]}), .init(2'b00), .state({trees[211], lumberyards[211]}));
acre acre_4_12 (.clk(clk), .en(en), .top_left({trees[161], lumberyards[161]}), .top({trees[162], lumberyards[162]}), .top_right({trees[163], lumberyards[163]}), .left({trees[211], lumberyards[211]}), .right({trees[213], lumberyards[213]}), .bottom_left({trees[261], lumberyards[261]}), .bottom({trees[262], lumberyards[262]}), .bottom_right({trees[263], lumberyards[263]}), .init(2'b00), .state({trees[212], lumberyards[212]}));
acre acre_4_13 (.clk(clk), .en(en), .top_left({trees[162], lumberyards[162]}), .top({trees[163], lumberyards[163]}), .top_right({trees[164], lumberyards[164]}), .left({trees[212], lumberyards[212]}), .right({trees[214], lumberyards[214]}), .bottom_left({trees[262], lumberyards[262]}), .bottom({trees[263], lumberyards[263]}), .bottom_right({trees[264], lumberyards[264]}), .init(2'b00), .state({trees[213], lumberyards[213]}));
acre acre_4_14 (.clk(clk), .en(en), .top_left({trees[163], lumberyards[163]}), .top({trees[164], lumberyards[164]}), .top_right({trees[165], lumberyards[165]}), .left({trees[213], lumberyards[213]}), .right({trees[215], lumberyards[215]}), .bottom_left({trees[263], lumberyards[263]}), .bottom({trees[264], lumberyards[264]}), .bottom_right({trees[265], lumberyards[265]}), .init(2'b00), .state({trees[214], lumberyards[214]}));
acre acre_4_15 (.clk(clk), .en(en), .top_left({trees[164], lumberyards[164]}), .top({trees[165], lumberyards[165]}), .top_right({trees[166], lumberyards[166]}), .left({trees[214], lumberyards[214]}), .right({trees[216], lumberyards[216]}), .bottom_left({trees[264], lumberyards[264]}), .bottom({trees[265], lumberyards[265]}), .bottom_right({trees[266], lumberyards[266]}), .init(2'b00), .state({trees[215], lumberyards[215]}));
acre acre_4_16 (.clk(clk), .en(en), .top_left({trees[165], lumberyards[165]}), .top({trees[166], lumberyards[166]}), .top_right({trees[167], lumberyards[167]}), .left({trees[215], lumberyards[215]}), .right({trees[217], lumberyards[217]}), .bottom_left({trees[265], lumberyards[265]}), .bottom({trees[266], lumberyards[266]}), .bottom_right({trees[267], lumberyards[267]}), .init(2'b10), .state({trees[216], lumberyards[216]}));
acre acre_4_17 (.clk(clk), .en(en), .top_left({trees[166], lumberyards[166]}), .top({trees[167], lumberyards[167]}), .top_right({trees[168], lumberyards[168]}), .left({trees[216], lumberyards[216]}), .right({trees[218], lumberyards[218]}), .bottom_left({trees[266], lumberyards[266]}), .bottom({trees[267], lumberyards[267]}), .bottom_right({trees[268], lumberyards[268]}), .init(2'b00), .state({trees[217], lumberyards[217]}));
acre acre_4_18 (.clk(clk), .en(en), .top_left({trees[167], lumberyards[167]}), .top({trees[168], lumberyards[168]}), .top_right({trees[169], lumberyards[169]}), .left({trees[217], lumberyards[217]}), .right({trees[219], lumberyards[219]}), .bottom_left({trees[267], lumberyards[267]}), .bottom({trees[268], lumberyards[268]}), .bottom_right({trees[269], lumberyards[269]}), .init(2'b00), .state({trees[218], lumberyards[218]}));
acre acre_4_19 (.clk(clk), .en(en), .top_left({trees[168], lumberyards[168]}), .top({trees[169], lumberyards[169]}), .top_right({trees[170], lumberyards[170]}), .left({trees[218], lumberyards[218]}), .right({trees[220], lumberyards[220]}), .bottom_left({trees[268], lumberyards[268]}), .bottom({trees[269], lumberyards[269]}), .bottom_right({trees[270], lumberyards[270]}), .init(2'b00), .state({trees[219], lumberyards[219]}));
acre acre_4_20 (.clk(clk), .en(en), .top_left({trees[169], lumberyards[169]}), .top({trees[170], lumberyards[170]}), .top_right({trees[171], lumberyards[171]}), .left({trees[219], lumberyards[219]}), .right({trees[221], lumberyards[221]}), .bottom_left({trees[269], lumberyards[269]}), .bottom({trees[270], lumberyards[270]}), .bottom_right({trees[271], lumberyards[271]}), .init(2'b10), .state({trees[220], lumberyards[220]}));
acre acre_4_21 (.clk(clk), .en(en), .top_left({trees[170], lumberyards[170]}), .top({trees[171], lumberyards[171]}), .top_right({trees[172], lumberyards[172]}), .left({trees[220], lumberyards[220]}), .right({trees[222], lumberyards[222]}), .bottom_left({trees[270], lumberyards[270]}), .bottom({trees[271], lumberyards[271]}), .bottom_right({trees[272], lumberyards[272]}), .init(2'b10), .state({trees[221], lumberyards[221]}));
acre acre_4_22 (.clk(clk), .en(en), .top_left({trees[171], lumberyards[171]}), .top({trees[172], lumberyards[172]}), .top_right({trees[173], lumberyards[173]}), .left({trees[221], lumberyards[221]}), .right({trees[223], lumberyards[223]}), .bottom_left({trees[271], lumberyards[271]}), .bottom({trees[272], lumberyards[272]}), .bottom_right({trees[273], lumberyards[273]}), .init(2'b01), .state({trees[222], lumberyards[222]}));
acre acre_4_23 (.clk(clk), .en(en), .top_left({trees[172], lumberyards[172]}), .top({trees[173], lumberyards[173]}), .top_right({trees[174], lumberyards[174]}), .left({trees[222], lumberyards[222]}), .right({trees[224], lumberyards[224]}), .bottom_left({trees[272], lumberyards[272]}), .bottom({trees[273], lumberyards[273]}), .bottom_right({trees[274], lumberyards[274]}), .init(2'b00), .state({trees[223], lumberyards[223]}));
acre acre_4_24 (.clk(clk), .en(en), .top_left({trees[173], lumberyards[173]}), .top({trees[174], lumberyards[174]}), .top_right({trees[175], lumberyards[175]}), .left({trees[223], lumberyards[223]}), .right({trees[225], lumberyards[225]}), .bottom_left({trees[273], lumberyards[273]}), .bottom({trees[274], lumberyards[274]}), .bottom_right({trees[275], lumberyards[275]}), .init(2'b01), .state({trees[224], lumberyards[224]}));
acre acre_4_25 (.clk(clk), .en(en), .top_left({trees[174], lumberyards[174]}), .top({trees[175], lumberyards[175]}), .top_right({trees[176], lumberyards[176]}), .left({trees[224], lumberyards[224]}), .right({trees[226], lumberyards[226]}), .bottom_left({trees[274], lumberyards[274]}), .bottom({trees[275], lumberyards[275]}), .bottom_right({trees[276], lumberyards[276]}), .init(2'b00), .state({trees[225], lumberyards[225]}));
acre acre_4_26 (.clk(clk), .en(en), .top_left({trees[175], lumberyards[175]}), .top({trees[176], lumberyards[176]}), .top_right({trees[177], lumberyards[177]}), .left({trees[225], lumberyards[225]}), .right({trees[227], lumberyards[227]}), .bottom_left({trees[275], lumberyards[275]}), .bottom({trees[276], lumberyards[276]}), .bottom_right({trees[277], lumberyards[277]}), .init(2'b00), .state({trees[226], lumberyards[226]}));
acre acre_4_27 (.clk(clk), .en(en), .top_left({trees[176], lumberyards[176]}), .top({trees[177], lumberyards[177]}), .top_right({trees[178], lumberyards[178]}), .left({trees[226], lumberyards[226]}), .right({trees[228], lumberyards[228]}), .bottom_left({trees[276], lumberyards[276]}), .bottom({trees[277], lumberyards[277]}), .bottom_right({trees[278], lumberyards[278]}), .init(2'b01), .state({trees[227], lumberyards[227]}));
acre acre_4_28 (.clk(clk), .en(en), .top_left({trees[177], lumberyards[177]}), .top({trees[178], lumberyards[178]}), .top_right({trees[179], lumberyards[179]}), .left({trees[227], lumberyards[227]}), .right({trees[229], lumberyards[229]}), .bottom_left({trees[277], lumberyards[277]}), .bottom({trees[278], lumberyards[278]}), .bottom_right({trees[279], lumberyards[279]}), .init(2'b01), .state({trees[228], lumberyards[228]}));
acre acre_4_29 (.clk(clk), .en(en), .top_left({trees[178], lumberyards[178]}), .top({trees[179], lumberyards[179]}), .top_right({trees[180], lumberyards[180]}), .left({trees[228], lumberyards[228]}), .right({trees[230], lumberyards[230]}), .bottom_left({trees[278], lumberyards[278]}), .bottom({trees[279], lumberyards[279]}), .bottom_right({trees[280], lumberyards[280]}), .init(2'b01), .state({trees[229], lumberyards[229]}));
acre acre_4_30 (.clk(clk), .en(en), .top_left({trees[179], lumberyards[179]}), .top({trees[180], lumberyards[180]}), .top_right({trees[181], lumberyards[181]}), .left({trees[229], lumberyards[229]}), .right({trees[231], lumberyards[231]}), .bottom_left({trees[279], lumberyards[279]}), .bottom({trees[280], lumberyards[280]}), .bottom_right({trees[281], lumberyards[281]}), .init(2'b00), .state({trees[230], lumberyards[230]}));
acre acre_4_31 (.clk(clk), .en(en), .top_left({trees[180], lumberyards[180]}), .top({trees[181], lumberyards[181]}), .top_right({trees[182], lumberyards[182]}), .left({trees[230], lumberyards[230]}), .right({trees[232], lumberyards[232]}), .bottom_left({trees[280], lumberyards[280]}), .bottom({trees[281], lumberyards[281]}), .bottom_right({trees[282], lumberyards[282]}), .init(2'b00), .state({trees[231], lumberyards[231]}));
acre acre_4_32 (.clk(clk), .en(en), .top_left({trees[181], lumberyards[181]}), .top({trees[182], lumberyards[182]}), .top_right({trees[183], lumberyards[183]}), .left({trees[231], lumberyards[231]}), .right({trees[233], lumberyards[233]}), .bottom_left({trees[281], lumberyards[281]}), .bottom({trees[282], lumberyards[282]}), .bottom_right({trees[283], lumberyards[283]}), .init(2'b01), .state({trees[232], lumberyards[232]}));
acre acre_4_33 (.clk(clk), .en(en), .top_left({trees[182], lumberyards[182]}), .top({trees[183], lumberyards[183]}), .top_right({trees[184], lumberyards[184]}), .left({trees[232], lumberyards[232]}), .right({trees[234], lumberyards[234]}), .bottom_left({trees[282], lumberyards[282]}), .bottom({trees[283], lumberyards[283]}), .bottom_right({trees[284], lumberyards[284]}), .init(2'b00), .state({trees[233], lumberyards[233]}));
acre acre_4_34 (.clk(clk), .en(en), .top_left({trees[183], lumberyards[183]}), .top({trees[184], lumberyards[184]}), .top_right({trees[185], lumberyards[185]}), .left({trees[233], lumberyards[233]}), .right({trees[235], lumberyards[235]}), .bottom_left({trees[283], lumberyards[283]}), .bottom({trees[284], lumberyards[284]}), .bottom_right({trees[285], lumberyards[285]}), .init(2'b00), .state({trees[234], lumberyards[234]}));
acre acre_4_35 (.clk(clk), .en(en), .top_left({trees[184], lumberyards[184]}), .top({trees[185], lumberyards[185]}), .top_right({trees[186], lumberyards[186]}), .left({trees[234], lumberyards[234]}), .right({trees[236], lumberyards[236]}), .bottom_left({trees[284], lumberyards[284]}), .bottom({trees[285], lumberyards[285]}), .bottom_right({trees[286], lumberyards[286]}), .init(2'b01), .state({trees[235], lumberyards[235]}));
acre acre_4_36 (.clk(clk), .en(en), .top_left({trees[185], lumberyards[185]}), .top({trees[186], lumberyards[186]}), .top_right({trees[187], lumberyards[187]}), .left({trees[235], lumberyards[235]}), .right({trees[237], lumberyards[237]}), .bottom_left({trees[285], lumberyards[285]}), .bottom({trees[286], lumberyards[286]}), .bottom_right({trees[287], lumberyards[287]}), .init(2'b01), .state({trees[236], lumberyards[236]}));
acre acre_4_37 (.clk(clk), .en(en), .top_left({trees[186], lumberyards[186]}), .top({trees[187], lumberyards[187]}), .top_right({trees[188], lumberyards[188]}), .left({trees[236], lumberyards[236]}), .right({trees[238], lumberyards[238]}), .bottom_left({trees[286], lumberyards[286]}), .bottom({trees[287], lumberyards[287]}), .bottom_right({trees[288], lumberyards[288]}), .init(2'b00), .state({trees[237], lumberyards[237]}));
acre acre_4_38 (.clk(clk), .en(en), .top_left({trees[187], lumberyards[187]}), .top({trees[188], lumberyards[188]}), .top_right({trees[189], lumberyards[189]}), .left({trees[237], lumberyards[237]}), .right({trees[239], lumberyards[239]}), .bottom_left({trees[287], lumberyards[287]}), .bottom({trees[288], lumberyards[288]}), .bottom_right({trees[289], lumberyards[289]}), .init(2'b00), .state({trees[238], lumberyards[238]}));
acre acre_4_39 (.clk(clk), .en(en), .top_left({trees[188], lumberyards[188]}), .top({trees[189], lumberyards[189]}), .top_right({trees[190], lumberyards[190]}), .left({trees[238], lumberyards[238]}), .right({trees[240], lumberyards[240]}), .bottom_left({trees[288], lumberyards[288]}), .bottom({trees[289], lumberyards[289]}), .bottom_right({trees[290], lumberyards[290]}), .init(2'b01), .state({trees[239], lumberyards[239]}));
acre acre_4_40 (.clk(clk), .en(en), .top_left({trees[189], lumberyards[189]}), .top({trees[190], lumberyards[190]}), .top_right({trees[191], lumberyards[191]}), .left({trees[239], lumberyards[239]}), .right({trees[241], lumberyards[241]}), .bottom_left({trees[289], lumberyards[289]}), .bottom({trees[290], lumberyards[290]}), .bottom_right({trees[291], lumberyards[291]}), .init(2'b00), .state({trees[240], lumberyards[240]}));
acre acre_4_41 (.clk(clk), .en(en), .top_left({trees[190], lumberyards[190]}), .top({trees[191], lumberyards[191]}), .top_right({trees[192], lumberyards[192]}), .left({trees[240], lumberyards[240]}), .right({trees[242], lumberyards[242]}), .bottom_left({trees[290], lumberyards[290]}), .bottom({trees[291], lumberyards[291]}), .bottom_right({trees[292], lumberyards[292]}), .init(2'b10), .state({trees[241], lumberyards[241]}));
acre acre_4_42 (.clk(clk), .en(en), .top_left({trees[191], lumberyards[191]}), .top({trees[192], lumberyards[192]}), .top_right({trees[193], lumberyards[193]}), .left({trees[241], lumberyards[241]}), .right({trees[243], lumberyards[243]}), .bottom_left({trees[291], lumberyards[291]}), .bottom({trees[292], lumberyards[292]}), .bottom_right({trees[293], lumberyards[293]}), .init(2'b10), .state({trees[242], lumberyards[242]}));
acre acre_4_43 (.clk(clk), .en(en), .top_left({trees[192], lumberyards[192]}), .top({trees[193], lumberyards[193]}), .top_right({trees[194], lumberyards[194]}), .left({trees[242], lumberyards[242]}), .right({trees[244], lumberyards[244]}), .bottom_left({trees[292], lumberyards[292]}), .bottom({trees[293], lumberyards[293]}), .bottom_right({trees[294], lumberyards[294]}), .init(2'b00), .state({trees[243], lumberyards[243]}));
acre acre_4_44 (.clk(clk), .en(en), .top_left({trees[193], lumberyards[193]}), .top({trees[194], lumberyards[194]}), .top_right({trees[195], lumberyards[195]}), .left({trees[243], lumberyards[243]}), .right({trees[245], lumberyards[245]}), .bottom_left({trees[293], lumberyards[293]}), .bottom({trees[294], lumberyards[294]}), .bottom_right({trees[295], lumberyards[295]}), .init(2'b00), .state({trees[244], lumberyards[244]}));
acre acre_4_45 (.clk(clk), .en(en), .top_left({trees[194], lumberyards[194]}), .top({trees[195], lumberyards[195]}), .top_right({trees[196], lumberyards[196]}), .left({trees[244], lumberyards[244]}), .right({trees[246], lumberyards[246]}), .bottom_left({trees[294], lumberyards[294]}), .bottom({trees[295], lumberyards[295]}), .bottom_right({trees[296], lumberyards[296]}), .init(2'b00), .state({trees[245], lumberyards[245]}));
acre acre_4_46 (.clk(clk), .en(en), .top_left({trees[195], lumberyards[195]}), .top({trees[196], lumberyards[196]}), .top_right({trees[197], lumberyards[197]}), .left({trees[245], lumberyards[245]}), .right({trees[247], lumberyards[247]}), .bottom_left({trees[295], lumberyards[295]}), .bottom({trees[296], lumberyards[296]}), .bottom_right({trees[297], lumberyards[297]}), .init(2'b01), .state({trees[246], lumberyards[246]}));
acre acre_4_47 (.clk(clk), .en(en), .top_left({trees[196], lumberyards[196]}), .top({trees[197], lumberyards[197]}), .top_right({trees[198], lumberyards[198]}), .left({trees[246], lumberyards[246]}), .right({trees[248], lumberyards[248]}), .bottom_left({trees[296], lumberyards[296]}), .bottom({trees[297], lumberyards[297]}), .bottom_right({trees[298], lumberyards[298]}), .init(2'b10), .state({trees[247], lumberyards[247]}));
acre acre_4_48 (.clk(clk), .en(en), .top_left({trees[197], lumberyards[197]}), .top({trees[198], lumberyards[198]}), .top_right({trees[199], lumberyards[199]}), .left({trees[247], lumberyards[247]}), .right({trees[249], lumberyards[249]}), .bottom_left({trees[297], lumberyards[297]}), .bottom({trees[298], lumberyards[298]}), .bottom_right({trees[299], lumberyards[299]}), .init(2'b01), .state({trees[248], lumberyards[248]}));
acre acre_4_49 (.clk(clk), .en(en), .top_left({trees[198], lumberyards[198]}), .top({trees[199], lumberyards[199]}), .top_right(2'b0), .left({trees[248], lumberyards[248]}), .right(2'b0), .bottom_left({trees[298], lumberyards[298]}), .bottom({trees[299], lumberyards[299]}), .bottom_right(2'b0), .init(2'b00), .state({trees[249], lumberyards[249]}));
acre acre_5_0 (.clk(clk), .en(en), .top_left(2'b0), .top({trees[200], lumberyards[200]}), .top_right({trees[201], lumberyards[201]}), .left(2'b0), .right({trees[251], lumberyards[251]}), .bottom_left(2'b0), .bottom({trees[300], lumberyards[300]}), .bottom_right({trees[301], lumberyards[301]}), .init(2'b00), .state({trees[250], lumberyards[250]}));
acre acre_5_1 (.clk(clk), .en(en), .top_left({trees[200], lumberyards[200]}), .top({trees[201], lumberyards[201]}), .top_right({trees[202], lumberyards[202]}), .left({trees[250], lumberyards[250]}), .right({trees[252], lumberyards[252]}), .bottom_left({trees[300], lumberyards[300]}), .bottom({trees[301], lumberyards[301]}), .bottom_right({trees[302], lumberyards[302]}), .init(2'b10), .state({trees[251], lumberyards[251]}));
acre acre_5_2 (.clk(clk), .en(en), .top_left({trees[201], lumberyards[201]}), .top({trees[202], lumberyards[202]}), .top_right({trees[203], lumberyards[203]}), .left({trees[251], lumberyards[251]}), .right({trees[253], lumberyards[253]}), .bottom_left({trees[301], lumberyards[301]}), .bottom({trees[302], lumberyards[302]}), .bottom_right({trees[303], lumberyards[303]}), .init(2'b10), .state({trees[252], lumberyards[252]}));
acre acre_5_3 (.clk(clk), .en(en), .top_left({trees[202], lumberyards[202]}), .top({trees[203], lumberyards[203]}), .top_right({trees[204], lumberyards[204]}), .left({trees[252], lumberyards[252]}), .right({trees[254], lumberyards[254]}), .bottom_left({trees[302], lumberyards[302]}), .bottom({trees[303], lumberyards[303]}), .bottom_right({trees[304], lumberyards[304]}), .init(2'b00), .state({trees[253], lumberyards[253]}));
acre acre_5_4 (.clk(clk), .en(en), .top_left({trees[203], lumberyards[203]}), .top({trees[204], lumberyards[204]}), .top_right({trees[205], lumberyards[205]}), .left({trees[253], lumberyards[253]}), .right({trees[255], lumberyards[255]}), .bottom_left({trees[303], lumberyards[303]}), .bottom({trees[304], lumberyards[304]}), .bottom_right({trees[305], lumberyards[305]}), .init(2'b00), .state({trees[254], lumberyards[254]}));
acre acre_5_5 (.clk(clk), .en(en), .top_left({trees[204], lumberyards[204]}), .top({trees[205], lumberyards[205]}), .top_right({trees[206], lumberyards[206]}), .left({trees[254], lumberyards[254]}), .right({trees[256], lumberyards[256]}), .bottom_left({trees[304], lumberyards[304]}), .bottom({trees[305], lumberyards[305]}), .bottom_right({trees[306], lumberyards[306]}), .init(2'b10), .state({trees[255], lumberyards[255]}));
acre acre_5_6 (.clk(clk), .en(en), .top_left({trees[205], lumberyards[205]}), .top({trees[206], lumberyards[206]}), .top_right({trees[207], lumberyards[207]}), .left({trees[255], lumberyards[255]}), .right({trees[257], lumberyards[257]}), .bottom_left({trees[305], lumberyards[305]}), .bottom({trees[306], lumberyards[306]}), .bottom_right({trees[307], lumberyards[307]}), .init(2'b00), .state({trees[256], lumberyards[256]}));
acre acre_5_7 (.clk(clk), .en(en), .top_left({trees[206], lumberyards[206]}), .top({trees[207], lumberyards[207]}), .top_right({trees[208], lumberyards[208]}), .left({trees[256], lumberyards[256]}), .right({trees[258], lumberyards[258]}), .bottom_left({trees[306], lumberyards[306]}), .bottom({trees[307], lumberyards[307]}), .bottom_right({trees[308], lumberyards[308]}), .init(2'b00), .state({trees[257], lumberyards[257]}));
acre acre_5_8 (.clk(clk), .en(en), .top_left({trees[207], lumberyards[207]}), .top({trees[208], lumberyards[208]}), .top_right({trees[209], lumberyards[209]}), .left({trees[257], lumberyards[257]}), .right({trees[259], lumberyards[259]}), .bottom_left({trees[307], lumberyards[307]}), .bottom({trees[308], lumberyards[308]}), .bottom_right({trees[309], lumberyards[309]}), .init(2'b00), .state({trees[258], lumberyards[258]}));
acre acre_5_9 (.clk(clk), .en(en), .top_left({trees[208], lumberyards[208]}), .top({trees[209], lumberyards[209]}), .top_right({trees[210], lumberyards[210]}), .left({trees[258], lumberyards[258]}), .right({trees[260], lumberyards[260]}), .bottom_left({trees[308], lumberyards[308]}), .bottom({trees[309], lumberyards[309]}), .bottom_right({trees[310], lumberyards[310]}), .init(2'b10), .state({trees[259], lumberyards[259]}));
acre acre_5_10 (.clk(clk), .en(en), .top_left({trees[209], lumberyards[209]}), .top({trees[210], lumberyards[210]}), .top_right({trees[211], lumberyards[211]}), .left({trees[259], lumberyards[259]}), .right({trees[261], lumberyards[261]}), .bottom_left({trees[309], lumberyards[309]}), .bottom({trees[310], lumberyards[310]}), .bottom_right({trees[311], lumberyards[311]}), .init(2'b10), .state({trees[260], lumberyards[260]}));
acre acre_5_11 (.clk(clk), .en(en), .top_left({trees[210], lumberyards[210]}), .top({trees[211], lumberyards[211]}), .top_right({trees[212], lumberyards[212]}), .left({trees[260], lumberyards[260]}), .right({trees[262], lumberyards[262]}), .bottom_left({trees[310], lumberyards[310]}), .bottom({trees[311], lumberyards[311]}), .bottom_right({trees[312], lumberyards[312]}), .init(2'b00), .state({trees[261], lumberyards[261]}));
acre acre_5_12 (.clk(clk), .en(en), .top_left({trees[211], lumberyards[211]}), .top({trees[212], lumberyards[212]}), .top_right({trees[213], lumberyards[213]}), .left({trees[261], lumberyards[261]}), .right({trees[263], lumberyards[263]}), .bottom_left({trees[311], lumberyards[311]}), .bottom({trees[312], lumberyards[312]}), .bottom_right({trees[313], lumberyards[313]}), .init(2'b00), .state({trees[262], lumberyards[262]}));
acre acre_5_13 (.clk(clk), .en(en), .top_left({trees[212], lumberyards[212]}), .top({trees[213], lumberyards[213]}), .top_right({trees[214], lumberyards[214]}), .left({trees[262], lumberyards[262]}), .right({trees[264], lumberyards[264]}), .bottom_left({trees[312], lumberyards[312]}), .bottom({trees[313], lumberyards[313]}), .bottom_right({trees[314], lumberyards[314]}), .init(2'b01), .state({trees[263], lumberyards[263]}));
acre acre_5_14 (.clk(clk), .en(en), .top_left({trees[213], lumberyards[213]}), .top({trees[214], lumberyards[214]}), .top_right({trees[215], lumberyards[215]}), .left({trees[263], lumberyards[263]}), .right({trees[265], lumberyards[265]}), .bottom_left({trees[313], lumberyards[313]}), .bottom({trees[314], lumberyards[314]}), .bottom_right({trees[315], lumberyards[315]}), .init(2'b00), .state({trees[264], lumberyards[264]}));
acre acre_5_15 (.clk(clk), .en(en), .top_left({trees[214], lumberyards[214]}), .top({trees[215], lumberyards[215]}), .top_right({trees[216], lumberyards[216]}), .left({trees[264], lumberyards[264]}), .right({trees[266], lumberyards[266]}), .bottom_left({trees[314], lumberyards[314]}), .bottom({trees[315], lumberyards[315]}), .bottom_right({trees[316], lumberyards[316]}), .init(2'b00), .state({trees[265], lumberyards[265]}));
acre acre_5_16 (.clk(clk), .en(en), .top_left({trees[215], lumberyards[215]}), .top({trees[216], lumberyards[216]}), .top_right({trees[217], lumberyards[217]}), .left({trees[265], lumberyards[265]}), .right({trees[267], lumberyards[267]}), .bottom_left({trees[315], lumberyards[315]}), .bottom({trees[316], lumberyards[316]}), .bottom_right({trees[317], lumberyards[317]}), .init(2'b00), .state({trees[266], lumberyards[266]}));
acre acre_5_17 (.clk(clk), .en(en), .top_left({trees[216], lumberyards[216]}), .top({trees[217], lumberyards[217]}), .top_right({trees[218], lumberyards[218]}), .left({trees[266], lumberyards[266]}), .right({trees[268], lumberyards[268]}), .bottom_left({trees[316], lumberyards[316]}), .bottom({trees[317], lumberyards[317]}), .bottom_right({trees[318], lumberyards[318]}), .init(2'b00), .state({trees[267], lumberyards[267]}));
acre acre_5_18 (.clk(clk), .en(en), .top_left({trees[217], lumberyards[217]}), .top({trees[218], lumberyards[218]}), .top_right({trees[219], lumberyards[219]}), .left({trees[267], lumberyards[267]}), .right({trees[269], lumberyards[269]}), .bottom_left({trees[317], lumberyards[317]}), .bottom({trees[318], lumberyards[318]}), .bottom_right({trees[319], lumberyards[319]}), .init(2'b00), .state({trees[268], lumberyards[268]}));
acre acre_5_19 (.clk(clk), .en(en), .top_left({trees[218], lumberyards[218]}), .top({trees[219], lumberyards[219]}), .top_right({trees[220], lumberyards[220]}), .left({trees[268], lumberyards[268]}), .right({trees[270], lumberyards[270]}), .bottom_left({trees[318], lumberyards[318]}), .bottom({trees[319], lumberyards[319]}), .bottom_right({trees[320], lumberyards[320]}), .init(2'b00), .state({trees[269], lumberyards[269]}));
acre acre_5_20 (.clk(clk), .en(en), .top_left({trees[219], lumberyards[219]}), .top({trees[220], lumberyards[220]}), .top_right({trees[221], lumberyards[221]}), .left({trees[269], lumberyards[269]}), .right({trees[271], lumberyards[271]}), .bottom_left({trees[319], lumberyards[319]}), .bottom({trees[320], lumberyards[320]}), .bottom_right({trees[321], lumberyards[321]}), .init(2'b01), .state({trees[270], lumberyards[270]}));
acre acre_5_21 (.clk(clk), .en(en), .top_left({trees[220], lumberyards[220]}), .top({trees[221], lumberyards[221]}), .top_right({trees[222], lumberyards[222]}), .left({trees[270], lumberyards[270]}), .right({trees[272], lumberyards[272]}), .bottom_left({trees[320], lumberyards[320]}), .bottom({trees[321], lumberyards[321]}), .bottom_right({trees[322], lumberyards[322]}), .init(2'b00), .state({trees[271], lumberyards[271]}));
acre acre_5_22 (.clk(clk), .en(en), .top_left({trees[221], lumberyards[221]}), .top({trees[222], lumberyards[222]}), .top_right({trees[223], lumberyards[223]}), .left({trees[271], lumberyards[271]}), .right({trees[273], lumberyards[273]}), .bottom_left({trees[321], lumberyards[321]}), .bottom({trees[322], lumberyards[322]}), .bottom_right({trees[323], lumberyards[323]}), .init(2'b01), .state({trees[272], lumberyards[272]}));
acre acre_5_23 (.clk(clk), .en(en), .top_left({trees[222], lumberyards[222]}), .top({trees[223], lumberyards[223]}), .top_right({trees[224], lumberyards[224]}), .left({trees[272], lumberyards[272]}), .right({trees[274], lumberyards[274]}), .bottom_left({trees[322], lumberyards[322]}), .bottom({trees[323], lumberyards[323]}), .bottom_right({trees[324], lumberyards[324]}), .init(2'b00), .state({trees[273], lumberyards[273]}));
acre acre_5_24 (.clk(clk), .en(en), .top_left({trees[223], lumberyards[223]}), .top({trees[224], lumberyards[224]}), .top_right({trees[225], lumberyards[225]}), .left({trees[273], lumberyards[273]}), .right({trees[275], lumberyards[275]}), .bottom_left({trees[323], lumberyards[323]}), .bottom({trees[324], lumberyards[324]}), .bottom_right({trees[325], lumberyards[325]}), .init(2'b00), .state({trees[274], lumberyards[274]}));
acre acre_5_25 (.clk(clk), .en(en), .top_left({trees[224], lumberyards[224]}), .top({trees[225], lumberyards[225]}), .top_right({trees[226], lumberyards[226]}), .left({trees[274], lumberyards[274]}), .right({trees[276], lumberyards[276]}), .bottom_left({trees[324], lumberyards[324]}), .bottom({trees[325], lumberyards[325]}), .bottom_right({trees[326], lumberyards[326]}), .init(2'b00), .state({trees[275], lumberyards[275]}));
acre acre_5_26 (.clk(clk), .en(en), .top_left({trees[225], lumberyards[225]}), .top({trees[226], lumberyards[226]}), .top_right({trees[227], lumberyards[227]}), .left({trees[275], lumberyards[275]}), .right({trees[277], lumberyards[277]}), .bottom_left({trees[325], lumberyards[325]}), .bottom({trees[326], lumberyards[326]}), .bottom_right({trees[327], lumberyards[327]}), .init(2'b00), .state({trees[276], lumberyards[276]}));
acre acre_5_27 (.clk(clk), .en(en), .top_left({trees[226], lumberyards[226]}), .top({trees[227], lumberyards[227]}), .top_right({trees[228], lumberyards[228]}), .left({trees[276], lumberyards[276]}), .right({trees[278], lumberyards[278]}), .bottom_left({trees[326], lumberyards[326]}), .bottom({trees[327], lumberyards[327]}), .bottom_right({trees[328], lumberyards[328]}), .init(2'b00), .state({trees[277], lumberyards[277]}));
acre acre_5_28 (.clk(clk), .en(en), .top_left({trees[227], lumberyards[227]}), .top({trees[228], lumberyards[228]}), .top_right({trees[229], lumberyards[229]}), .left({trees[277], lumberyards[277]}), .right({trees[279], lumberyards[279]}), .bottom_left({trees[327], lumberyards[327]}), .bottom({trees[328], lumberyards[328]}), .bottom_right({trees[329], lumberyards[329]}), .init(2'b00), .state({trees[278], lumberyards[278]}));
acre acre_5_29 (.clk(clk), .en(en), .top_left({trees[228], lumberyards[228]}), .top({trees[229], lumberyards[229]}), .top_right({trees[230], lumberyards[230]}), .left({trees[278], lumberyards[278]}), .right({trees[280], lumberyards[280]}), .bottom_left({trees[328], lumberyards[328]}), .bottom({trees[329], lumberyards[329]}), .bottom_right({trees[330], lumberyards[330]}), .init(2'b10), .state({trees[279], lumberyards[279]}));
acre acre_5_30 (.clk(clk), .en(en), .top_left({trees[229], lumberyards[229]}), .top({trees[230], lumberyards[230]}), .top_right({trees[231], lumberyards[231]}), .left({trees[279], lumberyards[279]}), .right({trees[281], lumberyards[281]}), .bottom_left({trees[329], lumberyards[329]}), .bottom({trees[330], lumberyards[330]}), .bottom_right({trees[331], lumberyards[331]}), .init(2'b00), .state({trees[280], lumberyards[280]}));
acre acre_5_31 (.clk(clk), .en(en), .top_left({trees[230], lumberyards[230]}), .top({trees[231], lumberyards[231]}), .top_right({trees[232], lumberyards[232]}), .left({trees[280], lumberyards[280]}), .right({trees[282], lumberyards[282]}), .bottom_left({trees[330], lumberyards[330]}), .bottom({trees[331], lumberyards[331]}), .bottom_right({trees[332], lumberyards[332]}), .init(2'b01), .state({trees[281], lumberyards[281]}));
acre acre_5_32 (.clk(clk), .en(en), .top_left({trees[231], lumberyards[231]}), .top({trees[232], lumberyards[232]}), .top_right({trees[233], lumberyards[233]}), .left({trees[281], lumberyards[281]}), .right({trees[283], lumberyards[283]}), .bottom_left({trees[331], lumberyards[331]}), .bottom({trees[332], lumberyards[332]}), .bottom_right({trees[333], lumberyards[333]}), .init(2'b00), .state({trees[282], lumberyards[282]}));
acre acre_5_33 (.clk(clk), .en(en), .top_left({trees[232], lumberyards[232]}), .top({trees[233], lumberyards[233]}), .top_right({trees[234], lumberyards[234]}), .left({trees[282], lumberyards[282]}), .right({trees[284], lumberyards[284]}), .bottom_left({trees[332], lumberyards[332]}), .bottom({trees[333], lumberyards[333]}), .bottom_right({trees[334], lumberyards[334]}), .init(2'b00), .state({trees[283], lumberyards[283]}));
acre acre_5_34 (.clk(clk), .en(en), .top_left({trees[233], lumberyards[233]}), .top({trees[234], lumberyards[234]}), .top_right({trees[235], lumberyards[235]}), .left({trees[283], lumberyards[283]}), .right({trees[285], lumberyards[285]}), .bottom_left({trees[333], lumberyards[333]}), .bottom({trees[334], lumberyards[334]}), .bottom_right({trees[335], lumberyards[335]}), .init(2'b00), .state({trees[284], lumberyards[284]}));
acre acre_5_35 (.clk(clk), .en(en), .top_left({trees[234], lumberyards[234]}), .top({trees[235], lumberyards[235]}), .top_right({trees[236], lumberyards[236]}), .left({trees[284], lumberyards[284]}), .right({trees[286], lumberyards[286]}), .bottom_left({trees[334], lumberyards[334]}), .bottom({trees[335], lumberyards[335]}), .bottom_right({trees[336], lumberyards[336]}), .init(2'b00), .state({trees[285], lumberyards[285]}));
acre acre_5_36 (.clk(clk), .en(en), .top_left({trees[235], lumberyards[235]}), .top({trees[236], lumberyards[236]}), .top_right({trees[237], lumberyards[237]}), .left({trees[285], lumberyards[285]}), .right({trees[287], lumberyards[287]}), .bottom_left({trees[335], lumberyards[335]}), .bottom({trees[336], lumberyards[336]}), .bottom_right({trees[337], lumberyards[337]}), .init(2'b10), .state({trees[286], lumberyards[286]}));
acre acre_5_37 (.clk(clk), .en(en), .top_left({trees[236], lumberyards[236]}), .top({trees[237], lumberyards[237]}), .top_right({trees[238], lumberyards[238]}), .left({trees[286], lumberyards[286]}), .right({trees[288], lumberyards[288]}), .bottom_left({trees[336], lumberyards[336]}), .bottom({trees[337], lumberyards[337]}), .bottom_right({trees[338], lumberyards[338]}), .init(2'b00), .state({trees[287], lumberyards[287]}));
acre acre_5_38 (.clk(clk), .en(en), .top_left({trees[237], lumberyards[237]}), .top({trees[238], lumberyards[238]}), .top_right({trees[239], lumberyards[239]}), .left({trees[287], lumberyards[287]}), .right({trees[289], lumberyards[289]}), .bottom_left({trees[337], lumberyards[337]}), .bottom({trees[338], lumberyards[338]}), .bottom_right({trees[339], lumberyards[339]}), .init(2'b01), .state({trees[288], lumberyards[288]}));
acre acre_5_39 (.clk(clk), .en(en), .top_left({trees[238], lumberyards[238]}), .top({trees[239], lumberyards[239]}), .top_right({trees[240], lumberyards[240]}), .left({trees[288], lumberyards[288]}), .right({trees[290], lumberyards[290]}), .bottom_left({trees[338], lumberyards[338]}), .bottom({trees[339], lumberyards[339]}), .bottom_right({trees[340], lumberyards[340]}), .init(2'b00), .state({trees[289], lumberyards[289]}));
acre acre_5_40 (.clk(clk), .en(en), .top_left({trees[239], lumberyards[239]}), .top({trees[240], lumberyards[240]}), .top_right({trees[241], lumberyards[241]}), .left({trees[289], lumberyards[289]}), .right({trees[291], lumberyards[291]}), .bottom_left({trees[339], lumberyards[339]}), .bottom({trees[340], lumberyards[340]}), .bottom_right({trees[341], lumberyards[341]}), .init(2'b00), .state({trees[290], lumberyards[290]}));
acre acre_5_41 (.clk(clk), .en(en), .top_left({trees[240], lumberyards[240]}), .top({trees[241], lumberyards[241]}), .top_right({trees[242], lumberyards[242]}), .left({trees[290], lumberyards[290]}), .right({trees[292], lumberyards[292]}), .bottom_left({trees[340], lumberyards[340]}), .bottom({trees[341], lumberyards[341]}), .bottom_right({trees[342], lumberyards[342]}), .init(2'b10), .state({trees[291], lumberyards[291]}));
acre acre_5_42 (.clk(clk), .en(en), .top_left({trees[241], lumberyards[241]}), .top({trees[242], lumberyards[242]}), .top_right({trees[243], lumberyards[243]}), .left({trees[291], lumberyards[291]}), .right({trees[293], lumberyards[293]}), .bottom_left({trees[341], lumberyards[341]}), .bottom({trees[342], lumberyards[342]}), .bottom_right({trees[343], lumberyards[343]}), .init(2'b00), .state({trees[292], lumberyards[292]}));
acre acre_5_43 (.clk(clk), .en(en), .top_left({trees[242], lumberyards[242]}), .top({trees[243], lumberyards[243]}), .top_right({trees[244], lumberyards[244]}), .left({trees[292], lumberyards[292]}), .right({trees[294], lumberyards[294]}), .bottom_left({trees[342], lumberyards[342]}), .bottom({trees[343], lumberyards[343]}), .bottom_right({trees[344], lumberyards[344]}), .init(2'b10), .state({trees[293], lumberyards[293]}));
acre acre_5_44 (.clk(clk), .en(en), .top_left({trees[243], lumberyards[243]}), .top({trees[244], lumberyards[244]}), .top_right({trees[245], lumberyards[245]}), .left({trees[293], lumberyards[293]}), .right({trees[295], lumberyards[295]}), .bottom_left({trees[343], lumberyards[343]}), .bottom({trees[344], lumberyards[344]}), .bottom_right({trees[345], lumberyards[345]}), .init(2'b00), .state({trees[294], lumberyards[294]}));
acre acre_5_45 (.clk(clk), .en(en), .top_left({trees[244], lumberyards[244]}), .top({trees[245], lumberyards[245]}), .top_right({trees[246], lumberyards[246]}), .left({trees[294], lumberyards[294]}), .right({trees[296], lumberyards[296]}), .bottom_left({trees[344], lumberyards[344]}), .bottom({trees[345], lumberyards[345]}), .bottom_right({trees[346], lumberyards[346]}), .init(2'b00), .state({trees[295], lumberyards[295]}));
acre acre_5_46 (.clk(clk), .en(en), .top_left({trees[245], lumberyards[245]}), .top({trees[246], lumberyards[246]}), .top_right({trees[247], lumberyards[247]}), .left({trees[295], lumberyards[295]}), .right({trees[297], lumberyards[297]}), .bottom_left({trees[345], lumberyards[345]}), .bottom({trees[346], lumberyards[346]}), .bottom_right({trees[347], lumberyards[347]}), .init(2'b10), .state({trees[296], lumberyards[296]}));
acre acre_5_47 (.clk(clk), .en(en), .top_left({trees[246], lumberyards[246]}), .top({trees[247], lumberyards[247]}), .top_right({trees[248], lumberyards[248]}), .left({trees[296], lumberyards[296]}), .right({trees[298], lumberyards[298]}), .bottom_left({trees[346], lumberyards[346]}), .bottom({trees[347], lumberyards[347]}), .bottom_right({trees[348], lumberyards[348]}), .init(2'b01), .state({trees[297], lumberyards[297]}));
acre acre_5_48 (.clk(clk), .en(en), .top_left({trees[247], lumberyards[247]}), .top({trees[248], lumberyards[248]}), .top_right({trees[249], lumberyards[249]}), .left({trees[297], lumberyards[297]}), .right({trees[299], lumberyards[299]}), .bottom_left({trees[347], lumberyards[347]}), .bottom({trees[348], lumberyards[348]}), .bottom_right({trees[349], lumberyards[349]}), .init(2'b00), .state({trees[298], lumberyards[298]}));
acre acre_5_49 (.clk(clk), .en(en), .top_left({trees[248], lumberyards[248]}), .top({trees[249], lumberyards[249]}), .top_right(2'b0), .left({trees[298], lumberyards[298]}), .right(2'b0), .bottom_left({trees[348], lumberyards[348]}), .bottom({trees[349], lumberyards[349]}), .bottom_right(2'b0), .init(2'b00), .state({trees[299], lumberyards[299]}));
acre acre_6_0 (.clk(clk), .en(en), .top_left(2'b0), .top({trees[250], lumberyards[250]}), .top_right({trees[251], lumberyards[251]}), .left(2'b0), .right({trees[301], lumberyards[301]}), .bottom_left(2'b0), .bottom({trees[350], lumberyards[350]}), .bottom_right({trees[351], lumberyards[351]}), .init(2'b00), .state({trees[300], lumberyards[300]}));
acre acre_6_1 (.clk(clk), .en(en), .top_left({trees[250], lumberyards[250]}), .top({trees[251], lumberyards[251]}), .top_right({trees[252], lumberyards[252]}), .left({trees[300], lumberyards[300]}), .right({trees[302], lumberyards[302]}), .bottom_left({trees[350], lumberyards[350]}), .bottom({trees[351], lumberyards[351]}), .bottom_right({trees[352], lumberyards[352]}), .init(2'b10), .state({trees[301], lumberyards[301]}));
acre acre_6_2 (.clk(clk), .en(en), .top_left({trees[251], lumberyards[251]}), .top({trees[252], lumberyards[252]}), .top_right({trees[253], lumberyards[253]}), .left({trees[301], lumberyards[301]}), .right({trees[303], lumberyards[303]}), .bottom_left({trees[351], lumberyards[351]}), .bottom({trees[352], lumberyards[352]}), .bottom_right({trees[353], lumberyards[353]}), .init(2'b00), .state({trees[302], lumberyards[302]}));
acre acre_6_3 (.clk(clk), .en(en), .top_left({trees[252], lumberyards[252]}), .top({trees[253], lumberyards[253]}), .top_right({trees[254], lumberyards[254]}), .left({trees[302], lumberyards[302]}), .right({trees[304], lumberyards[304]}), .bottom_left({trees[352], lumberyards[352]}), .bottom({trees[353], lumberyards[353]}), .bottom_right({trees[354], lumberyards[354]}), .init(2'b00), .state({trees[303], lumberyards[303]}));
acre acre_6_4 (.clk(clk), .en(en), .top_left({trees[253], lumberyards[253]}), .top({trees[254], lumberyards[254]}), .top_right({trees[255], lumberyards[255]}), .left({trees[303], lumberyards[303]}), .right({trees[305], lumberyards[305]}), .bottom_left({trees[353], lumberyards[353]}), .bottom({trees[354], lumberyards[354]}), .bottom_right({trees[355], lumberyards[355]}), .init(2'b00), .state({trees[304], lumberyards[304]}));
acre acre_6_5 (.clk(clk), .en(en), .top_left({trees[254], lumberyards[254]}), .top({trees[255], lumberyards[255]}), .top_right({trees[256], lumberyards[256]}), .left({trees[304], lumberyards[304]}), .right({trees[306], lumberyards[306]}), .bottom_left({trees[354], lumberyards[354]}), .bottom({trees[355], lumberyards[355]}), .bottom_right({trees[356], lumberyards[356]}), .init(2'b00), .state({trees[305], lumberyards[305]}));
acre acre_6_6 (.clk(clk), .en(en), .top_left({trees[255], lumberyards[255]}), .top({trees[256], lumberyards[256]}), .top_right({trees[257], lumberyards[257]}), .left({trees[305], lumberyards[305]}), .right({trees[307], lumberyards[307]}), .bottom_left({trees[355], lumberyards[355]}), .bottom({trees[356], lumberyards[356]}), .bottom_right({trees[357], lumberyards[357]}), .init(2'b00), .state({trees[306], lumberyards[306]}));
acre acre_6_7 (.clk(clk), .en(en), .top_left({trees[256], lumberyards[256]}), .top({trees[257], lumberyards[257]}), .top_right({trees[258], lumberyards[258]}), .left({trees[306], lumberyards[306]}), .right({trees[308], lumberyards[308]}), .bottom_left({trees[356], lumberyards[356]}), .bottom({trees[357], lumberyards[357]}), .bottom_right({trees[358], lumberyards[358]}), .init(2'b01), .state({trees[307], lumberyards[307]}));
acre acre_6_8 (.clk(clk), .en(en), .top_left({trees[257], lumberyards[257]}), .top({trees[258], lumberyards[258]}), .top_right({trees[259], lumberyards[259]}), .left({trees[307], lumberyards[307]}), .right({trees[309], lumberyards[309]}), .bottom_left({trees[357], lumberyards[357]}), .bottom({trees[358], lumberyards[358]}), .bottom_right({trees[359], lumberyards[359]}), .init(2'b10), .state({trees[308], lumberyards[308]}));
acre acre_6_9 (.clk(clk), .en(en), .top_left({trees[258], lumberyards[258]}), .top({trees[259], lumberyards[259]}), .top_right({trees[260], lumberyards[260]}), .left({trees[308], lumberyards[308]}), .right({trees[310], lumberyards[310]}), .bottom_left({trees[358], lumberyards[358]}), .bottom({trees[359], lumberyards[359]}), .bottom_right({trees[360], lumberyards[360]}), .init(2'b10), .state({trees[309], lumberyards[309]}));
acre acre_6_10 (.clk(clk), .en(en), .top_left({trees[259], lumberyards[259]}), .top({trees[260], lumberyards[260]}), .top_right({trees[261], lumberyards[261]}), .left({trees[309], lumberyards[309]}), .right({trees[311], lumberyards[311]}), .bottom_left({trees[359], lumberyards[359]}), .bottom({trees[360], lumberyards[360]}), .bottom_right({trees[361], lumberyards[361]}), .init(2'b00), .state({trees[310], lumberyards[310]}));
acre acre_6_11 (.clk(clk), .en(en), .top_left({trees[260], lumberyards[260]}), .top({trees[261], lumberyards[261]}), .top_right({trees[262], lumberyards[262]}), .left({trees[310], lumberyards[310]}), .right({trees[312], lumberyards[312]}), .bottom_left({trees[360], lumberyards[360]}), .bottom({trees[361], lumberyards[361]}), .bottom_right({trees[362], lumberyards[362]}), .init(2'b00), .state({trees[311], lumberyards[311]}));
acre acre_6_12 (.clk(clk), .en(en), .top_left({trees[261], lumberyards[261]}), .top({trees[262], lumberyards[262]}), .top_right({trees[263], lumberyards[263]}), .left({trees[311], lumberyards[311]}), .right({trees[313], lumberyards[313]}), .bottom_left({trees[361], lumberyards[361]}), .bottom({trees[362], lumberyards[362]}), .bottom_right({trees[363], lumberyards[363]}), .init(2'b00), .state({trees[312], lumberyards[312]}));
acre acre_6_13 (.clk(clk), .en(en), .top_left({trees[262], lumberyards[262]}), .top({trees[263], lumberyards[263]}), .top_right({trees[264], lumberyards[264]}), .left({trees[312], lumberyards[312]}), .right({trees[314], lumberyards[314]}), .bottom_left({trees[362], lumberyards[362]}), .bottom({trees[363], lumberyards[363]}), .bottom_right({trees[364], lumberyards[364]}), .init(2'b00), .state({trees[313], lumberyards[313]}));
acre acre_6_14 (.clk(clk), .en(en), .top_left({trees[263], lumberyards[263]}), .top({trees[264], lumberyards[264]}), .top_right({trees[265], lumberyards[265]}), .left({trees[313], lumberyards[313]}), .right({trees[315], lumberyards[315]}), .bottom_left({trees[363], lumberyards[363]}), .bottom({trees[364], lumberyards[364]}), .bottom_right({trees[365], lumberyards[365]}), .init(2'b00), .state({trees[314], lumberyards[314]}));
acre acre_6_15 (.clk(clk), .en(en), .top_left({trees[264], lumberyards[264]}), .top({trees[265], lumberyards[265]}), .top_right({trees[266], lumberyards[266]}), .left({trees[314], lumberyards[314]}), .right({trees[316], lumberyards[316]}), .bottom_left({trees[364], lumberyards[364]}), .bottom({trees[365], lumberyards[365]}), .bottom_right({trees[366], lumberyards[366]}), .init(2'b10), .state({trees[315], lumberyards[315]}));
acre acre_6_16 (.clk(clk), .en(en), .top_left({trees[265], lumberyards[265]}), .top({trees[266], lumberyards[266]}), .top_right({trees[267], lumberyards[267]}), .left({trees[315], lumberyards[315]}), .right({trees[317], lumberyards[317]}), .bottom_left({trees[365], lumberyards[365]}), .bottom({trees[366], lumberyards[366]}), .bottom_right({trees[367], lumberyards[367]}), .init(2'b01), .state({trees[316], lumberyards[316]}));
acre acre_6_17 (.clk(clk), .en(en), .top_left({trees[266], lumberyards[266]}), .top({trees[267], lumberyards[267]}), .top_right({trees[268], lumberyards[268]}), .left({trees[316], lumberyards[316]}), .right({trees[318], lumberyards[318]}), .bottom_left({trees[366], lumberyards[366]}), .bottom({trees[367], lumberyards[367]}), .bottom_right({trees[368], lumberyards[368]}), .init(2'b00), .state({trees[317], lumberyards[317]}));
acre acre_6_18 (.clk(clk), .en(en), .top_left({trees[267], lumberyards[267]}), .top({trees[268], lumberyards[268]}), .top_right({trees[269], lumberyards[269]}), .left({trees[317], lumberyards[317]}), .right({trees[319], lumberyards[319]}), .bottom_left({trees[367], lumberyards[367]}), .bottom({trees[368], lumberyards[368]}), .bottom_right({trees[369], lumberyards[369]}), .init(2'b01), .state({trees[318], lumberyards[318]}));
acre acre_6_19 (.clk(clk), .en(en), .top_left({trees[268], lumberyards[268]}), .top({trees[269], lumberyards[269]}), .top_right({trees[270], lumberyards[270]}), .left({trees[318], lumberyards[318]}), .right({trees[320], lumberyards[320]}), .bottom_left({trees[368], lumberyards[368]}), .bottom({trees[369], lumberyards[369]}), .bottom_right({trees[370], lumberyards[370]}), .init(2'b01), .state({trees[319], lumberyards[319]}));
acre acre_6_20 (.clk(clk), .en(en), .top_left({trees[269], lumberyards[269]}), .top({trees[270], lumberyards[270]}), .top_right({trees[271], lumberyards[271]}), .left({trees[319], lumberyards[319]}), .right({trees[321], lumberyards[321]}), .bottom_left({trees[369], lumberyards[369]}), .bottom({trees[370], lumberyards[370]}), .bottom_right({trees[371], lumberyards[371]}), .init(2'b01), .state({trees[320], lumberyards[320]}));
acre acre_6_21 (.clk(clk), .en(en), .top_left({trees[270], lumberyards[270]}), .top({trees[271], lumberyards[271]}), .top_right({trees[272], lumberyards[272]}), .left({trees[320], lumberyards[320]}), .right({trees[322], lumberyards[322]}), .bottom_left({trees[370], lumberyards[370]}), .bottom({trees[371], lumberyards[371]}), .bottom_right({trees[372], lumberyards[372]}), .init(2'b00), .state({trees[321], lumberyards[321]}));
acre acre_6_22 (.clk(clk), .en(en), .top_left({trees[271], lumberyards[271]}), .top({trees[272], lumberyards[272]}), .top_right({trees[273], lumberyards[273]}), .left({trees[321], lumberyards[321]}), .right({trees[323], lumberyards[323]}), .bottom_left({trees[371], lumberyards[371]}), .bottom({trees[372], lumberyards[372]}), .bottom_right({trees[373], lumberyards[373]}), .init(2'b00), .state({trees[322], lumberyards[322]}));
acre acre_6_23 (.clk(clk), .en(en), .top_left({trees[272], lumberyards[272]}), .top({trees[273], lumberyards[273]}), .top_right({trees[274], lumberyards[274]}), .left({trees[322], lumberyards[322]}), .right({trees[324], lumberyards[324]}), .bottom_left({trees[372], lumberyards[372]}), .bottom({trees[373], lumberyards[373]}), .bottom_right({trees[374], lumberyards[374]}), .init(2'b00), .state({trees[323], lumberyards[323]}));
acre acre_6_24 (.clk(clk), .en(en), .top_left({trees[273], lumberyards[273]}), .top({trees[274], lumberyards[274]}), .top_right({trees[275], lumberyards[275]}), .left({trees[323], lumberyards[323]}), .right({trees[325], lumberyards[325]}), .bottom_left({trees[373], lumberyards[373]}), .bottom({trees[374], lumberyards[374]}), .bottom_right({trees[375], lumberyards[375]}), .init(2'b00), .state({trees[324], lumberyards[324]}));
acre acre_6_25 (.clk(clk), .en(en), .top_left({trees[274], lumberyards[274]}), .top({trees[275], lumberyards[275]}), .top_right({trees[276], lumberyards[276]}), .left({trees[324], lumberyards[324]}), .right({trees[326], lumberyards[326]}), .bottom_left({trees[374], lumberyards[374]}), .bottom({trees[375], lumberyards[375]}), .bottom_right({trees[376], lumberyards[376]}), .init(2'b01), .state({trees[325], lumberyards[325]}));
acre acre_6_26 (.clk(clk), .en(en), .top_left({trees[275], lumberyards[275]}), .top({trees[276], lumberyards[276]}), .top_right({trees[277], lumberyards[277]}), .left({trees[325], lumberyards[325]}), .right({trees[327], lumberyards[327]}), .bottom_left({trees[375], lumberyards[375]}), .bottom({trees[376], lumberyards[376]}), .bottom_right({trees[377], lumberyards[377]}), .init(2'b00), .state({trees[326], lumberyards[326]}));
acre acre_6_27 (.clk(clk), .en(en), .top_left({trees[276], lumberyards[276]}), .top({trees[277], lumberyards[277]}), .top_right({trees[278], lumberyards[278]}), .left({trees[326], lumberyards[326]}), .right({trees[328], lumberyards[328]}), .bottom_left({trees[376], lumberyards[376]}), .bottom({trees[377], lumberyards[377]}), .bottom_right({trees[378], lumberyards[378]}), .init(2'b00), .state({trees[327], lumberyards[327]}));
acre acre_6_28 (.clk(clk), .en(en), .top_left({trees[277], lumberyards[277]}), .top({trees[278], lumberyards[278]}), .top_right({trees[279], lumberyards[279]}), .left({trees[327], lumberyards[327]}), .right({trees[329], lumberyards[329]}), .bottom_left({trees[377], lumberyards[377]}), .bottom({trees[378], lumberyards[378]}), .bottom_right({trees[379], lumberyards[379]}), .init(2'b01), .state({trees[328], lumberyards[328]}));
acre acre_6_29 (.clk(clk), .en(en), .top_left({trees[278], lumberyards[278]}), .top({trees[279], lumberyards[279]}), .top_right({trees[280], lumberyards[280]}), .left({trees[328], lumberyards[328]}), .right({trees[330], lumberyards[330]}), .bottom_left({trees[378], lumberyards[378]}), .bottom({trees[379], lumberyards[379]}), .bottom_right({trees[380], lumberyards[380]}), .init(2'b01), .state({trees[329], lumberyards[329]}));
acre acre_6_30 (.clk(clk), .en(en), .top_left({trees[279], lumberyards[279]}), .top({trees[280], lumberyards[280]}), .top_right({trees[281], lumberyards[281]}), .left({trees[329], lumberyards[329]}), .right({trees[331], lumberyards[331]}), .bottom_left({trees[379], lumberyards[379]}), .bottom({trees[380], lumberyards[380]}), .bottom_right({trees[381], lumberyards[381]}), .init(2'b00), .state({trees[330], lumberyards[330]}));
acre acre_6_31 (.clk(clk), .en(en), .top_left({trees[280], lumberyards[280]}), .top({trees[281], lumberyards[281]}), .top_right({trees[282], lumberyards[282]}), .left({trees[330], lumberyards[330]}), .right({trees[332], lumberyards[332]}), .bottom_left({trees[380], lumberyards[380]}), .bottom({trees[381], lumberyards[381]}), .bottom_right({trees[382], lumberyards[382]}), .init(2'b00), .state({trees[331], lumberyards[331]}));
acre acre_6_32 (.clk(clk), .en(en), .top_left({trees[281], lumberyards[281]}), .top({trees[282], lumberyards[282]}), .top_right({trees[283], lumberyards[283]}), .left({trees[331], lumberyards[331]}), .right({trees[333], lumberyards[333]}), .bottom_left({trees[381], lumberyards[381]}), .bottom({trees[382], lumberyards[382]}), .bottom_right({trees[383], lumberyards[383]}), .init(2'b01), .state({trees[332], lumberyards[332]}));
acre acre_6_33 (.clk(clk), .en(en), .top_left({trees[282], lumberyards[282]}), .top({trees[283], lumberyards[283]}), .top_right({trees[284], lumberyards[284]}), .left({trees[332], lumberyards[332]}), .right({trees[334], lumberyards[334]}), .bottom_left({trees[382], lumberyards[382]}), .bottom({trees[383], lumberyards[383]}), .bottom_right({trees[384], lumberyards[384]}), .init(2'b10), .state({trees[333], lumberyards[333]}));
acre acre_6_34 (.clk(clk), .en(en), .top_left({trees[283], lumberyards[283]}), .top({trees[284], lumberyards[284]}), .top_right({trees[285], lumberyards[285]}), .left({trees[333], lumberyards[333]}), .right({trees[335], lumberyards[335]}), .bottom_left({trees[383], lumberyards[383]}), .bottom({trees[384], lumberyards[384]}), .bottom_right({trees[385], lumberyards[385]}), .init(2'b01), .state({trees[334], lumberyards[334]}));
acre acre_6_35 (.clk(clk), .en(en), .top_left({trees[284], lumberyards[284]}), .top({trees[285], lumberyards[285]}), .top_right({trees[286], lumberyards[286]}), .left({trees[334], lumberyards[334]}), .right({trees[336], lumberyards[336]}), .bottom_left({trees[384], lumberyards[384]}), .bottom({trees[385], lumberyards[385]}), .bottom_right({trees[386], lumberyards[386]}), .init(2'b00), .state({trees[335], lumberyards[335]}));
acre acre_6_36 (.clk(clk), .en(en), .top_left({trees[285], lumberyards[285]}), .top({trees[286], lumberyards[286]}), .top_right({trees[287], lumberyards[287]}), .left({trees[335], lumberyards[335]}), .right({trees[337], lumberyards[337]}), .bottom_left({trees[385], lumberyards[385]}), .bottom({trees[386], lumberyards[386]}), .bottom_right({trees[387], lumberyards[387]}), .init(2'b00), .state({trees[336], lumberyards[336]}));
acre acre_6_37 (.clk(clk), .en(en), .top_left({trees[286], lumberyards[286]}), .top({trees[287], lumberyards[287]}), .top_right({trees[288], lumberyards[288]}), .left({trees[336], lumberyards[336]}), .right({trees[338], lumberyards[338]}), .bottom_left({trees[386], lumberyards[386]}), .bottom({trees[387], lumberyards[387]}), .bottom_right({trees[388], lumberyards[388]}), .init(2'b00), .state({trees[337], lumberyards[337]}));
acre acre_6_38 (.clk(clk), .en(en), .top_left({trees[287], lumberyards[287]}), .top({trees[288], lumberyards[288]}), .top_right({trees[289], lumberyards[289]}), .left({trees[337], lumberyards[337]}), .right({trees[339], lumberyards[339]}), .bottom_left({trees[387], lumberyards[387]}), .bottom({trees[388], lumberyards[388]}), .bottom_right({trees[389], lumberyards[389]}), .init(2'b10), .state({trees[338], lumberyards[338]}));
acre acre_6_39 (.clk(clk), .en(en), .top_left({trees[288], lumberyards[288]}), .top({trees[289], lumberyards[289]}), .top_right({trees[290], lumberyards[290]}), .left({trees[338], lumberyards[338]}), .right({trees[340], lumberyards[340]}), .bottom_left({trees[388], lumberyards[388]}), .bottom({trees[389], lumberyards[389]}), .bottom_right({trees[390], lumberyards[390]}), .init(2'b01), .state({trees[339], lumberyards[339]}));
acre acre_6_40 (.clk(clk), .en(en), .top_left({trees[289], lumberyards[289]}), .top({trees[290], lumberyards[290]}), .top_right({trees[291], lumberyards[291]}), .left({trees[339], lumberyards[339]}), .right({trees[341], lumberyards[341]}), .bottom_left({trees[389], lumberyards[389]}), .bottom({trees[390], lumberyards[390]}), .bottom_right({trees[391], lumberyards[391]}), .init(2'b01), .state({trees[340], lumberyards[340]}));
acre acre_6_41 (.clk(clk), .en(en), .top_left({trees[290], lumberyards[290]}), .top({trees[291], lumberyards[291]}), .top_right({trees[292], lumberyards[292]}), .left({trees[340], lumberyards[340]}), .right({trees[342], lumberyards[342]}), .bottom_left({trees[390], lumberyards[390]}), .bottom({trees[391], lumberyards[391]}), .bottom_right({trees[392], lumberyards[392]}), .init(2'b00), .state({trees[341], lumberyards[341]}));
acre acre_6_42 (.clk(clk), .en(en), .top_left({trees[291], lumberyards[291]}), .top({trees[292], lumberyards[292]}), .top_right({trees[293], lumberyards[293]}), .left({trees[341], lumberyards[341]}), .right({trees[343], lumberyards[343]}), .bottom_left({trees[391], lumberyards[391]}), .bottom({trees[392], lumberyards[392]}), .bottom_right({trees[393], lumberyards[393]}), .init(2'b00), .state({trees[342], lumberyards[342]}));
acre acre_6_43 (.clk(clk), .en(en), .top_left({trees[292], lumberyards[292]}), .top({trees[293], lumberyards[293]}), .top_right({trees[294], lumberyards[294]}), .left({trees[342], lumberyards[342]}), .right({trees[344], lumberyards[344]}), .bottom_left({trees[392], lumberyards[392]}), .bottom({trees[393], lumberyards[393]}), .bottom_right({trees[394], lumberyards[394]}), .init(2'b00), .state({trees[343], lumberyards[343]}));
acre acre_6_44 (.clk(clk), .en(en), .top_left({trees[293], lumberyards[293]}), .top({trees[294], lumberyards[294]}), .top_right({trees[295], lumberyards[295]}), .left({trees[343], lumberyards[343]}), .right({trees[345], lumberyards[345]}), .bottom_left({trees[393], lumberyards[393]}), .bottom({trees[394], lumberyards[394]}), .bottom_right({trees[395], lumberyards[395]}), .init(2'b00), .state({trees[344], lumberyards[344]}));
acre acre_6_45 (.clk(clk), .en(en), .top_left({trees[294], lumberyards[294]}), .top({trees[295], lumberyards[295]}), .top_right({trees[296], lumberyards[296]}), .left({trees[344], lumberyards[344]}), .right({trees[346], lumberyards[346]}), .bottom_left({trees[394], lumberyards[394]}), .bottom({trees[395], lumberyards[395]}), .bottom_right({trees[396], lumberyards[396]}), .init(2'b01), .state({trees[345], lumberyards[345]}));
acre acre_6_46 (.clk(clk), .en(en), .top_left({trees[295], lumberyards[295]}), .top({trees[296], lumberyards[296]}), .top_right({trees[297], lumberyards[297]}), .left({trees[345], lumberyards[345]}), .right({trees[347], lumberyards[347]}), .bottom_left({trees[395], lumberyards[395]}), .bottom({trees[396], lumberyards[396]}), .bottom_right({trees[397], lumberyards[397]}), .init(2'b10), .state({trees[346], lumberyards[346]}));
acre acre_6_47 (.clk(clk), .en(en), .top_left({trees[296], lumberyards[296]}), .top({trees[297], lumberyards[297]}), .top_right({trees[298], lumberyards[298]}), .left({trees[346], lumberyards[346]}), .right({trees[348], lumberyards[348]}), .bottom_left({trees[396], lumberyards[396]}), .bottom({trees[397], lumberyards[397]}), .bottom_right({trees[398], lumberyards[398]}), .init(2'b00), .state({trees[347], lumberyards[347]}));
acre acre_6_48 (.clk(clk), .en(en), .top_left({trees[297], lumberyards[297]}), .top({trees[298], lumberyards[298]}), .top_right({trees[299], lumberyards[299]}), .left({trees[347], lumberyards[347]}), .right({trees[349], lumberyards[349]}), .bottom_left({trees[397], lumberyards[397]}), .bottom({trees[398], lumberyards[398]}), .bottom_right({trees[399], lumberyards[399]}), .init(2'b01), .state({trees[348], lumberyards[348]}));
acre acre_6_49 (.clk(clk), .en(en), .top_left({trees[298], lumberyards[298]}), .top({trees[299], lumberyards[299]}), .top_right(2'b0), .left({trees[348], lumberyards[348]}), .right(2'b0), .bottom_left({trees[398], lumberyards[398]}), .bottom({trees[399], lumberyards[399]}), .bottom_right(2'b0), .init(2'b00), .state({trees[349], lumberyards[349]}));
acre acre_7_0 (.clk(clk), .en(en), .top_left(2'b0), .top({trees[300], lumberyards[300]}), .top_right({trees[301], lumberyards[301]}), .left(2'b0), .right({trees[351], lumberyards[351]}), .bottom_left(2'b0), .bottom({trees[400], lumberyards[400]}), .bottom_right({trees[401], lumberyards[401]}), .init(2'b00), .state({trees[350], lumberyards[350]}));
acre acre_7_1 (.clk(clk), .en(en), .top_left({trees[300], lumberyards[300]}), .top({trees[301], lumberyards[301]}), .top_right({trees[302], lumberyards[302]}), .left({trees[350], lumberyards[350]}), .right({trees[352], lumberyards[352]}), .bottom_left({trees[400], lumberyards[400]}), .bottom({trees[401], lumberyards[401]}), .bottom_right({trees[402], lumberyards[402]}), .init(2'b10), .state({trees[351], lumberyards[351]}));
acre acre_7_2 (.clk(clk), .en(en), .top_left({trees[301], lumberyards[301]}), .top({trees[302], lumberyards[302]}), .top_right({trees[303], lumberyards[303]}), .left({trees[351], lumberyards[351]}), .right({trees[353], lumberyards[353]}), .bottom_left({trees[401], lumberyards[401]}), .bottom({trees[402], lumberyards[402]}), .bottom_right({trees[403], lumberyards[403]}), .init(2'b01), .state({trees[352], lumberyards[352]}));
acre acre_7_3 (.clk(clk), .en(en), .top_left({trees[302], lumberyards[302]}), .top({trees[303], lumberyards[303]}), .top_right({trees[304], lumberyards[304]}), .left({trees[352], lumberyards[352]}), .right({trees[354], lumberyards[354]}), .bottom_left({trees[402], lumberyards[402]}), .bottom({trees[403], lumberyards[403]}), .bottom_right({trees[404], lumberyards[404]}), .init(2'b00), .state({trees[353], lumberyards[353]}));
acre acre_7_4 (.clk(clk), .en(en), .top_left({trees[303], lumberyards[303]}), .top({trees[304], lumberyards[304]}), .top_right({trees[305], lumberyards[305]}), .left({trees[353], lumberyards[353]}), .right({trees[355], lumberyards[355]}), .bottom_left({trees[403], lumberyards[403]}), .bottom({trees[404], lumberyards[404]}), .bottom_right({trees[405], lumberyards[405]}), .init(2'b00), .state({trees[354], lumberyards[354]}));
acre acre_7_5 (.clk(clk), .en(en), .top_left({trees[304], lumberyards[304]}), .top({trees[305], lumberyards[305]}), .top_right({trees[306], lumberyards[306]}), .left({trees[354], lumberyards[354]}), .right({trees[356], lumberyards[356]}), .bottom_left({trees[404], lumberyards[404]}), .bottom({trees[405], lumberyards[405]}), .bottom_right({trees[406], lumberyards[406]}), .init(2'b00), .state({trees[355], lumberyards[355]}));
acre acre_7_6 (.clk(clk), .en(en), .top_left({trees[305], lumberyards[305]}), .top({trees[306], lumberyards[306]}), .top_right({trees[307], lumberyards[307]}), .left({trees[355], lumberyards[355]}), .right({trees[357], lumberyards[357]}), .bottom_left({trees[405], lumberyards[405]}), .bottom({trees[406], lumberyards[406]}), .bottom_right({trees[407], lumberyards[407]}), .init(2'b00), .state({trees[356], lumberyards[356]}));
acre acre_7_7 (.clk(clk), .en(en), .top_left({trees[306], lumberyards[306]}), .top({trees[307], lumberyards[307]}), .top_right({trees[308], lumberyards[308]}), .left({trees[356], lumberyards[356]}), .right({trees[358], lumberyards[358]}), .bottom_left({trees[406], lumberyards[406]}), .bottom({trees[407], lumberyards[407]}), .bottom_right({trees[408], lumberyards[408]}), .init(2'b00), .state({trees[357], lumberyards[357]}));
acre acre_7_8 (.clk(clk), .en(en), .top_left({trees[307], lumberyards[307]}), .top({trees[308], lumberyards[308]}), .top_right({trees[309], lumberyards[309]}), .left({trees[357], lumberyards[357]}), .right({trees[359], lumberyards[359]}), .bottom_left({trees[407], lumberyards[407]}), .bottom({trees[408], lumberyards[408]}), .bottom_right({trees[409], lumberyards[409]}), .init(2'b00), .state({trees[358], lumberyards[358]}));
acre acre_7_9 (.clk(clk), .en(en), .top_left({trees[308], lumberyards[308]}), .top({trees[309], lumberyards[309]}), .top_right({trees[310], lumberyards[310]}), .left({trees[358], lumberyards[358]}), .right({trees[360], lumberyards[360]}), .bottom_left({trees[408], lumberyards[408]}), .bottom({trees[409], lumberyards[409]}), .bottom_right({trees[410], lumberyards[410]}), .init(2'b10), .state({trees[359], lumberyards[359]}));
acre acre_7_10 (.clk(clk), .en(en), .top_left({trees[309], lumberyards[309]}), .top({trees[310], lumberyards[310]}), .top_right({trees[311], lumberyards[311]}), .left({trees[359], lumberyards[359]}), .right({trees[361], lumberyards[361]}), .bottom_left({trees[409], lumberyards[409]}), .bottom({trees[410], lumberyards[410]}), .bottom_right({trees[411], lumberyards[411]}), .init(2'b10), .state({trees[360], lumberyards[360]}));
acre acre_7_11 (.clk(clk), .en(en), .top_left({trees[310], lumberyards[310]}), .top({trees[311], lumberyards[311]}), .top_right({trees[312], lumberyards[312]}), .left({trees[360], lumberyards[360]}), .right({trees[362], lumberyards[362]}), .bottom_left({trees[410], lumberyards[410]}), .bottom({trees[411], lumberyards[411]}), .bottom_right({trees[412], lumberyards[412]}), .init(2'b00), .state({trees[361], lumberyards[361]}));
acre acre_7_12 (.clk(clk), .en(en), .top_left({trees[311], lumberyards[311]}), .top({trees[312], lumberyards[312]}), .top_right({trees[313], lumberyards[313]}), .left({trees[361], lumberyards[361]}), .right({trees[363], lumberyards[363]}), .bottom_left({trees[411], lumberyards[411]}), .bottom({trees[412], lumberyards[412]}), .bottom_right({trees[413], lumberyards[413]}), .init(2'b00), .state({trees[362], lumberyards[362]}));
acre acre_7_13 (.clk(clk), .en(en), .top_left({trees[312], lumberyards[312]}), .top({trees[313], lumberyards[313]}), .top_right({trees[314], lumberyards[314]}), .left({trees[362], lumberyards[362]}), .right({trees[364], lumberyards[364]}), .bottom_left({trees[412], lumberyards[412]}), .bottom({trees[413], lumberyards[413]}), .bottom_right({trees[414], lumberyards[414]}), .init(2'b00), .state({trees[363], lumberyards[363]}));
acre acre_7_14 (.clk(clk), .en(en), .top_left({trees[313], lumberyards[313]}), .top({trees[314], lumberyards[314]}), .top_right({trees[315], lumberyards[315]}), .left({trees[363], lumberyards[363]}), .right({trees[365], lumberyards[365]}), .bottom_left({trees[413], lumberyards[413]}), .bottom({trees[414], lumberyards[414]}), .bottom_right({trees[415], lumberyards[415]}), .init(2'b00), .state({trees[364], lumberyards[364]}));
acre acre_7_15 (.clk(clk), .en(en), .top_left({trees[314], lumberyards[314]}), .top({trees[315], lumberyards[315]}), .top_right({trees[316], lumberyards[316]}), .left({trees[364], lumberyards[364]}), .right({trees[366], lumberyards[366]}), .bottom_left({trees[414], lumberyards[414]}), .bottom({trees[415], lumberyards[415]}), .bottom_right({trees[416], lumberyards[416]}), .init(2'b10), .state({trees[365], lumberyards[365]}));
acre acre_7_16 (.clk(clk), .en(en), .top_left({trees[315], lumberyards[315]}), .top({trees[316], lumberyards[316]}), .top_right({trees[317], lumberyards[317]}), .left({trees[365], lumberyards[365]}), .right({trees[367], lumberyards[367]}), .bottom_left({trees[415], lumberyards[415]}), .bottom({trees[416], lumberyards[416]}), .bottom_right({trees[417], lumberyards[417]}), .init(2'b01), .state({trees[366], lumberyards[366]}));
acre acre_7_17 (.clk(clk), .en(en), .top_left({trees[316], lumberyards[316]}), .top({trees[317], lumberyards[317]}), .top_right({trees[318], lumberyards[318]}), .left({trees[366], lumberyards[366]}), .right({trees[368], lumberyards[368]}), .bottom_left({trees[416], lumberyards[416]}), .bottom({trees[417], lumberyards[417]}), .bottom_right({trees[418], lumberyards[418]}), .init(2'b00), .state({trees[367], lumberyards[367]}));
acre acre_7_18 (.clk(clk), .en(en), .top_left({trees[317], lumberyards[317]}), .top({trees[318], lumberyards[318]}), .top_right({trees[319], lumberyards[319]}), .left({trees[367], lumberyards[367]}), .right({trees[369], lumberyards[369]}), .bottom_left({trees[417], lumberyards[417]}), .bottom({trees[418], lumberyards[418]}), .bottom_right({trees[419], lumberyards[419]}), .init(2'b00), .state({trees[368], lumberyards[368]}));
acre acre_7_19 (.clk(clk), .en(en), .top_left({trees[318], lumberyards[318]}), .top({trees[319], lumberyards[319]}), .top_right({trees[320], lumberyards[320]}), .left({trees[368], lumberyards[368]}), .right({trees[370], lumberyards[370]}), .bottom_left({trees[418], lumberyards[418]}), .bottom({trees[419], lumberyards[419]}), .bottom_right({trees[420], lumberyards[420]}), .init(2'b00), .state({trees[369], lumberyards[369]}));
acre acre_7_20 (.clk(clk), .en(en), .top_left({trees[319], lumberyards[319]}), .top({trees[320], lumberyards[320]}), .top_right({trees[321], lumberyards[321]}), .left({trees[369], lumberyards[369]}), .right({trees[371], lumberyards[371]}), .bottom_left({trees[419], lumberyards[419]}), .bottom({trees[420], lumberyards[420]}), .bottom_right({trees[421], lumberyards[421]}), .init(2'b01), .state({trees[370], lumberyards[370]}));
acre acre_7_21 (.clk(clk), .en(en), .top_left({trees[320], lumberyards[320]}), .top({trees[321], lumberyards[321]}), .top_right({trees[322], lumberyards[322]}), .left({trees[370], lumberyards[370]}), .right({trees[372], lumberyards[372]}), .bottom_left({trees[420], lumberyards[420]}), .bottom({trees[421], lumberyards[421]}), .bottom_right({trees[422], lumberyards[422]}), .init(2'b01), .state({trees[371], lumberyards[371]}));
acre acre_7_22 (.clk(clk), .en(en), .top_left({trees[321], lumberyards[321]}), .top({trees[322], lumberyards[322]}), .top_right({trees[323], lumberyards[323]}), .left({trees[371], lumberyards[371]}), .right({trees[373], lumberyards[373]}), .bottom_left({trees[421], lumberyards[421]}), .bottom({trees[422], lumberyards[422]}), .bottom_right({trees[423], lumberyards[423]}), .init(2'b00), .state({trees[372], lumberyards[372]}));
acre acre_7_23 (.clk(clk), .en(en), .top_left({trees[322], lumberyards[322]}), .top({trees[323], lumberyards[323]}), .top_right({trees[324], lumberyards[324]}), .left({trees[372], lumberyards[372]}), .right({trees[374], lumberyards[374]}), .bottom_left({trees[422], lumberyards[422]}), .bottom({trees[423], lumberyards[423]}), .bottom_right({trees[424], lumberyards[424]}), .init(2'b01), .state({trees[373], lumberyards[373]}));
acre acre_7_24 (.clk(clk), .en(en), .top_left({trees[323], lumberyards[323]}), .top({trees[324], lumberyards[324]}), .top_right({trees[325], lumberyards[325]}), .left({trees[373], lumberyards[373]}), .right({trees[375], lumberyards[375]}), .bottom_left({trees[423], lumberyards[423]}), .bottom({trees[424], lumberyards[424]}), .bottom_right({trees[425], lumberyards[425]}), .init(2'b00), .state({trees[374], lumberyards[374]}));
acre acre_7_25 (.clk(clk), .en(en), .top_left({trees[324], lumberyards[324]}), .top({trees[325], lumberyards[325]}), .top_right({trees[326], lumberyards[326]}), .left({trees[374], lumberyards[374]}), .right({trees[376], lumberyards[376]}), .bottom_left({trees[424], lumberyards[424]}), .bottom({trees[425], lumberyards[425]}), .bottom_right({trees[426], lumberyards[426]}), .init(2'b00), .state({trees[375], lumberyards[375]}));
acre acre_7_26 (.clk(clk), .en(en), .top_left({trees[325], lumberyards[325]}), .top({trees[326], lumberyards[326]}), .top_right({trees[327], lumberyards[327]}), .left({trees[375], lumberyards[375]}), .right({trees[377], lumberyards[377]}), .bottom_left({trees[425], lumberyards[425]}), .bottom({trees[426], lumberyards[426]}), .bottom_right({trees[427], lumberyards[427]}), .init(2'b00), .state({trees[376], lumberyards[376]}));
acre acre_7_27 (.clk(clk), .en(en), .top_left({trees[326], lumberyards[326]}), .top({trees[327], lumberyards[327]}), .top_right({trees[328], lumberyards[328]}), .left({trees[376], lumberyards[376]}), .right({trees[378], lumberyards[378]}), .bottom_left({trees[426], lumberyards[426]}), .bottom({trees[427], lumberyards[427]}), .bottom_right({trees[428], lumberyards[428]}), .init(2'b10), .state({trees[377], lumberyards[377]}));
acre acre_7_28 (.clk(clk), .en(en), .top_left({trees[327], lumberyards[327]}), .top({trees[328], lumberyards[328]}), .top_right({trees[329], lumberyards[329]}), .left({trees[377], lumberyards[377]}), .right({trees[379], lumberyards[379]}), .bottom_left({trees[427], lumberyards[427]}), .bottom({trees[428], lumberyards[428]}), .bottom_right({trees[429], lumberyards[429]}), .init(2'b00), .state({trees[378], lumberyards[378]}));
acre acre_7_29 (.clk(clk), .en(en), .top_left({trees[328], lumberyards[328]}), .top({trees[329], lumberyards[329]}), .top_right({trees[330], lumberyards[330]}), .left({trees[378], lumberyards[378]}), .right({trees[380], lumberyards[380]}), .bottom_left({trees[428], lumberyards[428]}), .bottom({trees[429], lumberyards[429]}), .bottom_right({trees[430], lumberyards[430]}), .init(2'b00), .state({trees[379], lumberyards[379]}));
acre acre_7_30 (.clk(clk), .en(en), .top_left({trees[329], lumberyards[329]}), .top({trees[330], lumberyards[330]}), .top_right({trees[331], lumberyards[331]}), .left({trees[379], lumberyards[379]}), .right({trees[381], lumberyards[381]}), .bottom_left({trees[429], lumberyards[429]}), .bottom({trees[430], lumberyards[430]}), .bottom_right({trees[431], lumberyards[431]}), .init(2'b00), .state({trees[380], lumberyards[380]}));
acre acre_7_31 (.clk(clk), .en(en), .top_left({trees[330], lumberyards[330]}), .top({trees[331], lumberyards[331]}), .top_right({trees[332], lumberyards[332]}), .left({trees[380], lumberyards[380]}), .right({trees[382], lumberyards[382]}), .bottom_left({trees[430], lumberyards[430]}), .bottom({trees[431], lumberyards[431]}), .bottom_right({trees[432], lumberyards[432]}), .init(2'b00), .state({trees[381], lumberyards[381]}));
acre acre_7_32 (.clk(clk), .en(en), .top_left({trees[331], lumberyards[331]}), .top({trees[332], lumberyards[332]}), .top_right({trees[333], lumberyards[333]}), .left({trees[381], lumberyards[381]}), .right({trees[383], lumberyards[383]}), .bottom_left({trees[431], lumberyards[431]}), .bottom({trees[432], lumberyards[432]}), .bottom_right({trees[433], lumberyards[433]}), .init(2'b10), .state({trees[382], lumberyards[382]}));
acre acre_7_33 (.clk(clk), .en(en), .top_left({trees[332], lumberyards[332]}), .top({trees[333], lumberyards[333]}), .top_right({trees[334], lumberyards[334]}), .left({trees[382], lumberyards[382]}), .right({trees[384], lumberyards[384]}), .bottom_left({trees[432], lumberyards[432]}), .bottom({trees[433], lumberyards[433]}), .bottom_right({trees[434], lumberyards[434]}), .init(2'b00), .state({trees[383], lumberyards[383]}));
acre acre_7_34 (.clk(clk), .en(en), .top_left({trees[333], lumberyards[333]}), .top({trees[334], lumberyards[334]}), .top_right({trees[335], lumberyards[335]}), .left({trees[383], lumberyards[383]}), .right({trees[385], lumberyards[385]}), .bottom_left({trees[433], lumberyards[433]}), .bottom({trees[434], lumberyards[434]}), .bottom_right({trees[435], lumberyards[435]}), .init(2'b01), .state({trees[384], lumberyards[384]}));
acre acre_7_35 (.clk(clk), .en(en), .top_left({trees[334], lumberyards[334]}), .top({trees[335], lumberyards[335]}), .top_right({trees[336], lumberyards[336]}), .left({trees[384], lumberyards[384]}), .right({trees[386], lumberyards[386]}), .bottom_left({trees[434], lumberyards[434]}), .bottom({trees[435], lumberyards[435]}), .bottom_right({trees[436], lumberyards[436]}), .init(2'b00), .state({trees[385], lumberyards[385]}));
acre acre_7_36 (.clk(clk), .en(en), .top_left({trees[335], lumberyards[335]}), .top({trees[336], lumberyards[336]}), .top_right({trees[337], lumberyards[337]}), .left({trees[385], lumberyards[385]}), .right({trees[387], lumberyards[387]}), .bottom_left({trees[435], lumberyards[435]}), .bottom({trees[436], lumberyards[436]}), .bottom_right({trees[437], lumberyards[437]}), .init(2'b00), .state({trees[386], lumberyards[386]}));
acre acre_7_37 (.clk(clk), .en(en), .top_left({trees[336], lumberyards[336]}), .top({trees[337], lumberyards[337]}), .top_right({trees[338], lumberyards[338]}), .left({trees[386], lumberyards[386]}), .right({trees[388], lumberyards[388]}), .bottom_left({trees[436], lumberyards[436]}), .bottom({trees[437], lumberyards[437]}), .bottom_right({trees[438], lumberyards[438]}), .init(2'b00), .state({trees[387], lumberyards[387]}));
acre acre_7_38 (.clk(clk), .en(en), .top_left({trees[337], lumberyards[337]}), .top({trees[338], lumberyards[338]}), .top_right({trees[339], lumberyards[339]}), .left({trees[387], lumberyards[387]}), .right({trees[389], lumberyards[389]}), .bottom_left({trees[437], lumberyards[437]}), .bottom({trees[438], lumberyards[438]}), .bottom_right({trees[439], lumberyards[439]}), .init(2'b00), .state({trees[388], lumberyards[388]}));
acre acre_7_39 (.clk(clk), .en(en), .top_left({trees[338], lumberyards[338]}), .top({trees[339], lumberyards[339]}), .top_right({trees[340], lumberyards[340]}), .left({trees[388], lumberyards[388]}), .right({trees[390], lumberyards[390]}), .bottom_left({trees[438], lumberyards[438]}), .bottom({trees[439], lumberyards[439]}), .bottom_right({trees[440], lumberyards[440]}), .init(2'b00), .state({trees[389], lumberyards[389]}));
acre acre_7_40 (.clk(clk), .en(en), .top_left({trees[339], lumberyards[339]}), .top({trees[340], lumberyards[340]}), .top_right({trees[341], lumberyards[341]}), .left({trees[389], lumberyards[389]}), .right({trees[391], lumberyards[391]}), .bottom_left({trees[439], lumberyards[439]}), .bottom({trees[440], lumberyards[440]}), .bottom_right({trees[441], lumberyards[441]}), .init(2'b00), .state({trees[390], lumberyards[390]}));
acre acre_7_41 (.clk(clk), .en(en), .top_left({trees[340], lumberyards[340]}), .top({trees[341], lumberyards[341]}), .top_right({trees[342], lumberyards[342]}), .left({trees[390], lumberyards[390]}), .right({trees[392], lumberyards[392]}), .bottom_left({trees[440], lumberyards[440]}), .bottom({trees[441], lumberyards[441]}), .bottom_right({trees[442], lumberyards[442]}), .init(2'b10), .state({trees[391], lumberyards[391]}));
acre acre_7_42 (.clk(clk), .en(en), .top_left({trees[341], lumberyards[341]}), .top({trees[342], lumberyards[342]}), .top_right({trees[343], lumberyards[343]}), .left({trees[391], lumberyards[391]}), .right({trees[393], lumberyards[393]}), .bottom_left({trees[441], lumberyards[441]}), .bottom({trees[442], lumberyards[442]}), .bottom_right({trees[443], lumberyards[443]}), .init(2'b00), .state({trees[392], lumberyards[392]}));
acre acre_7_43 (.clk(clk), .en(en), .top_left({trees[342], lumberyards[342]}), .top({trees[343], lumberyards[343]}), .top_right({trees[344], lumberyards[344]}), .left({trees[392], lumberyards[392]}), .right({trees[394], lumberyards[394]}), .bottom_left({trees[442], lumberyards[442]}), .bottom({trees[443], lumberyards[443]}), .bottom_right({trees[444], lumberyards[444]}), .init(2'b00), .state({trees[393], lumberyards[393]}));
acre acre_7_44 (.clk(clk), .en(en), .top_left({trees[343], lumberyards[343]}), .top({trees[344], lumberyards[344]}), .top_right({trees[345], lumberyards[345]}), .left({trees[393], lumberyards[393]}), .right({trees[395], lumberyards[395]}), .bottom_left({trees[443], lumberyards[443]}), .bottom({trees[444], lumberyards[444]}), .bottom_right({trees[445], lumberyards[445]}), .init(2'b00), .state({trees[394], lumberyards[394]}));
acre acre_7_45 (.clk(clk), .en(en), .top_left({trees[344], lumberyards[344]}), .top({trees[345], lumberyards[345]}), .top_right({trees[346], lumberyards[346]}), .left({trees[394], lumberyards[394]}), .right({trees[396], lumberyards[396]}), .bottom_left({trees[444], lumberyards[444]}), .bottom({trees[445], lumberyards[445]}), .bottom_right({trees[446], lumberyards[446]}), .init(2'b00), .state({trees[395], lumberyards[395]}));
acre acre_7_46 (.clk(clk), .en(en), .top_left({trees[345], lumberyards[345]}), .top({trees[346], lumberyards[346]}), .top_right({trees[347], lumberyards[347]}), .left({trees[395], lumberyards[395]}), .right({trees[397], lumberyards[397]}), .bottom_left({trees[445], lumberyards[445]}), .bottom({trees[446], lumberyards[446]}), .bottom_right({trees[447], lumberyards[447]}), .init(2'b00), .state({trees[396], lumberyards[396]}));
acre acre_7_47 (.clk(clk), .en(en), .top_left({trees[346], lumberyards[346]}), .top({trees[347], lumberyards[347]}), .top_right({trees[348], lumberyards[348]}), .left({trees[396], lumberyards[396]}), .right({trees[398], lumberyards[398]}), .bottom_left({trees[446], lumberyards[446]}), .bottom({trees[447], lumberyards[447]}), .bottom_right({trees[448], lumberyards[448]}), .init(2'b01), .state({trees[397], lumberyards[397]}));
acre acre_7_48 (.clk(clk), .en(en), .top_left({trees[347], lumberyards[347]}), .top({trees[348], lumberyards[348]}), .top_right({trees[349], lumberyards[349]}), .left({trees[397], lumberyards[397]}), .right({trees[399], lumberyards[399]}), .bottom_left({trees[447], lumberyards[447]}), .bottom({trees[448], lumberyards[448]}), .bottom_right({trees[449], lumberyards[449]}), .init(2'b00), .state({trees[398], lumberyards[398]}));
acre acre_7_49 (.clk(clk), .en(en), .top_left({trees[348], lumberyards[348]}), .top({trees[349], lumberyards[349]}), .top_right(2'b0), .left({trees[398], lumberyards[398]}), .right(2'b0), .bottom_left({trees[448], lumberyards[448]}), .bottom({trees[449], lumberyards[449]}), .bottom_right(2'b0), .init(2'b00), .state({trees[399], lumberyards[399]}));
acre acre_8_0 (.clk(clk), .en(en), .top_left(2'b0), .top({trees[350], lumberyards[350]}), .top_right({trees[351], lumberyards[351]}), .left(2'b0), .right({trees[401], lumberyards[401]}), .bottom_left(2'b0), .bottom({trees[450], lumberyards[450]}), .bottom_right({trees[451], lumberyards[451]}), .init(2'b01), .state({trees[400], lumberyards[400]}));
acre acre_8_1 (.clk(clk), .en(en), .top_left({trees[350], lumberyards[350]}), .top({trees[351], lumberyards[351]}), .top_right({trees[352], lumberyards[352]}), .left({trees[400], lumberyards[400]}), .right({trees[402], lumberyards[402]}), .bottom_left({trees[450], lumberyards[450]}), .bottom({trees[451], lumberyards[451]}), .bottom_right({trees[452], lumberyards[452]}), .init(2'b01), .state({trees[401], lumberyards[401]}));
acre acre_8_2 (.clk(clk), .en(en), .top_left({trees[351], lumberyards[351]}), .top({trees[352], lumberyards[352]}), .top_right({trees[353], lumberyards[353]}), .left({trees[401], lumberyards[401]}), .right({trees[403], lumberyards[403]}), .bottom_left({trees[451], lumberyards[451]}), .bottom({trees[452], lumberyards[452]}), .bottom_right({trees[453], lumberyards[453]}), .init(2'b00), .state({trees[402], lumberyards[402]}));
acre acre_8_3 (.clk(clk), .en(en), .top_left({trees[352], lumberyards[352]}), .top({trees[353], lumberyards[353]}), .top_right({trees[354], lumberyards[354]}), .left({trees[402], lumberyards[402]}), .right({trees[404], lumberyards[404]}), .bottom_left({trees[452], lumberyards[452]}), .bottom({trees[453], lumberyards[453]}), .bottom_right({trees[454], lumberyards[454]}), .init(2'b00), .state({trees[403], lumberyards[403]}));
acre acre_8_4 (.clk(clk), .en(en), .top_left({trees[353], lumberyards[353]}), .top({trees[354], lumberyards[354]}), .top_right({trees[355], lumberyards[355]}), .left({trees[403], lumberyards[403]}), .right({trees[405], lumberyards[405]}), .bottom_left({trees[453], lumberyards[453]}), .bottom({trees[454], lumberyards[454]}), .bottom_right({trees[455], lumberyards[455]}), .init(2'b10), .state({trees[404], lumberyards[404]}));
acre acre_8_5 (.clk(clk), .en(en), .top_left({trees[354], lumberyards[354]}), .top({trees[355], lumberyards[355]}), .top_right({trees[356], lumberyards[356]}), .left({trees[404], lumberyards[404]}), .right({trees[406], lumberyards[406]}), .bottom_left({trees[454], lumberyards[454]}), .bottom({trees[455], lumberyards[455]}), .bottom_right({trees[456], lumberyards[456]}), .init(2'b10), .state({trees[405], lumberyards[405]}));
acre acre_8_6 (.clk(clk), .en(en), .top_left({trees[355], lumberyards[355]}), .top({trees[356], lumberyards[356]}), .top_right({trees[357], lumberyards[357]}), .left({trees[405], lumberyards[405]}), .right({trees[407], lumberyards[407]}), .bottom_left({trees[455], lumberyards[455]}), .bottom({trees[456], lumberyards[456]}), .bottom_right({trees[457], lumberyards[457]}), .init(2'b00), .state({trees[406], lumberyards[406]}));
acre acre_8_7 (.clk(clk), .en(en), .top_left({trees[356], lumberyards[356]}), .top({trees[357], lumberyards[357]}), .top_right({trees[358], lumberyards[358]}), .left({trees[406], lumberyards[406]}), .right({trees[408], lumberyards[408]}), .bottom_left({trees[456], lumberyards[456]}), .bottom({trees[457], lumberyards[457]}), .bottom_right({trees[458], lumberyards[458]}), .init(2'b00), .state({trees[407], lumberyards[407]}));
acre acre_8_8 (.clk(clk), .en(en), .top_left({trees[357], lumberyards[357]}), .top({trees[358], lumberyards[358]}), .top_right({trees[359], lumberyards[359]}), .left({trees[407], lumberyards[407]}), .right({trees[409], lumberyards[409]}), .bottom_left({trees[457], lumberyards[457]}), .bottom({trees[458], lumberyards[458]}), .bottom_right({trees[459], lumberyards[459]}), .init(2'b01), .state({trees[408], lumberyards[408]}));
acre acre_8_9 (.clk(clk), .en(en), .top_left({trees[358], lumberyards[358]}), .top({trees[359], lumberyards[359]}), .top_right({trees[360], lumberyards[360]}), .left({trees[408], lumberyards[408]}), .right({trees[410], lumberyards[410]}), .bottom_left({trees[458], lumberyards[458]}), .bottom({trees[459], lumberyards[459]}), .bottom_right({trees[460], lumberyards[460]}), .init(2'b00), .state({trees[409], lumberyards[409]}));
acre acre_8_10 (.clk(clk), .en(en), .top_left({trees[359], lumberyards[359]}), .top({trees[360], lumberyards[360]}), .top_right({trees[361], lumberyards[361]}), .left({trees[409], lumberyards[409]}), .right({trees[411], lumberyards[411]}), .bottom_left({trees[459], lumberyards[459]}), .bottom({trees[460], lumberyards[460]}), .bottom_right({trees[461], lumberyards[461]}), .init(2'b00), .state({trees[410], lumberyards[410]}));
acre acre_8_11 (.clk(clk), .en(en), .top_left({trees[360], lumberyards[360]}), .top({trees[361], lumberyards[361]}), .top_right({trees[362], lumberyards[362]}), .left({trees[410], lumberyards[410]}), .right({trees[412], lumberyards[412]}), .bottom_left({trees[460], lumberyards[460]}), .bottom({trees[461], lumberyards[461]}), .bottom_right({trees[462], lumberyards[462]}), .init(2'b00), .state({trees[411], lumberyards[411]}));
acre acre_8_12 (.clk(clk), .en(en), .top_left({trees[361], lumberyards[361]}), .top({trees[362], lumberyards[362]}), .top_right({trees[363], lumberyards[363]}), .left({trees[411], lumberyards[411]}), .right({trees[413], lumberyards[413]}), .bottom_left({trees[461], lumberyards[461]}), .bottom({trees[462], lumberyards[462]}), .bottom_right({trees[463], lumberyards[463]}), .init(2'b01), .state({trees[412], lumberyards[412]}));
acre acre_8_13 (.clk(clk), .en(en), .top_left({trees[362], lumberyards[362]}), .top({trees[363], lumberyards[363]}), .top_right({trees[364], lumberyards[364]}), .left({trees[412], lumberyards[412]}), .right({trees[414], lumberyards[414]}), .bottom_left({trees[462], lumberyards[462]}), .bottom({trees[463], lumberyards[463]}), .bottom_right({trees[464], lumberyards[464]}), .init(2'b00), .state({trees[413], lumberyards[413]}));
acre acre_8_14 (.clk(clk), .en(en), .top_left({trees[363], lumberyards[363]}), .top({trees[364], lumberyards[364]}), .top_right({trees[365], lumberyards[365]}), .left({trees[413], lumberyards[413]}), .right({trees[415], lumberyards[415]}), .bottom_left({trees[463], lumberyards[463]}), .bottom({trees[464], lumberyards[464]}), .bottom_right({trees[465], lumberyards[465]}), .init(2'b00), .state({trees[414], lumberyards[414]}));
acre acre_8_15 (.clk(clk), .en(en), .top_left({trees[364], lumberyards[364]}), .top({trees[365], lumberyards[365]}), .top_right({trees[366], lumberyards[366]}), .left({trees[414], lumberyards[414]}), .right({trees[416], lumberyards[416]}), .bottom_left({trees[464], lumberyards[464]}), .bottom({trees[465], lumberyards[465]}), .bottom_right({trees[466], lumberyards[466]}), .init(2'b00), .state({trees[415], lumberyards[415]}));
acre acre_8_16 (.clk(clk), .en(en), .top_left({trees[365], lumberyards[365]}), .top({trees[366], lumberyards[366]}), .top_right({trees[367], lumberyards[367]}), .left({trees[415], lumberyards[415]}), .right({trees[417], lumberyards[417]}), .bottom_left({trees[465], lumberyards[465]}), .bottom({trees[466], lumberyards[466]}), .bottom_right({trees[467], lumberyards[467]}), .init(2'b00), .state({trees[416], lumberyards[416]}));
acre acre_8_17 (.clk(clk), .en(en), .top_left({trees[366], lumberyards[366]}), .top({trees[367], lumberyards[367]}), .top_right({trees[368], lumberyards[368]}), .left({trees[416], lumberyards[416]}), .right({trees[418], lumberyards[418]}), .bottom_left({trees[466], lumberyards[466]}), .bottom({trees[467], lumberyards[467]}), .bottom_right({trees[468], lumberyards[468]}), .init(2'b00), .state({trees[417], lumberyards[417]}));
acre acre_8_18 (.clk(clk), .en(en), .top_left({trees[367], lumberyards[367]}), .top({trees[368], lumberyards[368]}), .top_right({trees[369], lumberyards[369]}), .left({trees[417], lumberyards[417]}), .right({trees[419], lumberyards[419]}), .bottom_left({trees[467], lumberyards[467]}), .bottom({trees[468], lumberyards[468]}), .bottom_right({trees[469], lumberyards[469]}), .init(2'b00), .state({trees[418], lumberyards[418]}));
acre acre_8_19 (.clk(clk), .en(en), .top_left({trees[368], lumberyards[368]}), .top({trees[369], lumberyards[369]}), .top_right({trees[370], lumberyards[370]}), .left({trees[418], lumberyards[418]}), .right({trees[420], lumberyards[420]}), .bottom_left({trees[468], lumberyards[468]}), .bottom({trees[469], lumberyards[469]}), .bottom_right({trees[470], lumberyards[470]}), .init(2'b00), .state({trees[419], lumberyards[419]}));
acre acre_8_20 (.clk(clk), .en(en), .top_left({trees[369], lumberyards[369]}), .top({trees[370], lumberyards[370]}), .top_right({trees[371], lumberyards[371]}), .left({trees[419], lumberyards[419]}), .right({trees[421], lumberyards[421]}), .bottom_left({trees[469], lumberyards[469]}), .bottom({trees[470], lumberyards[470]}), .bottom_right({trees[471], lumberyards[471]}), .init(2'b00), .state({trees[420], lumberyards[420]}));
acre acre_8_21 (.clk(clk), .en(en), .top_left({trees[370], lumberyards[370]}), .top({trees[371], lumberyards[371]}), .top_right({trees[372], lumberyards[372]}), .left({trees[420], lumberyards[420]}), .right({trees[422], lumberyards[422]}), .bottom_left({trees[470], lumberyards[470]}), .bottom({trees[471], lumberyards[471]}), .bottom_right({trees[472], lumberyards[472]}), .init(2'b10), .state({trees[421], lumberyards[421]}));
acre acre_8_22 (.clk(clk), .en(en), .top_left({trees[371], lumberyards[371]}), .top({trees[372], lumberyards[372]}), .top_right({trees[373], lumberyards[373]}), .left({trees[421], lumberyards[421]}), .right({trees[423], lumberyards[423]}), .bottom_left({trees[471], lumberyards[471]}), .bottom({trees[472], lumberyards[472]}), .bottom_right({trees[473], lumberyards[473]}), .init(2'b00), .state({trees[422], lumberyards[422]}));
acre acre_8_23 (.clk(clk), .en(en), .top_left({trees[372], lumberyards[372]}), .top({trees[373], lumberyards[373]}), .top_right({trees[374], lumberyards[374]}), .left({trees[422], lumberyards[422]}), .right({trees[424], lumberyards[424]}), .bottom_left({trees[472], lumberyards[472]}), .bottom({trees[473], lumberyards[473]}), .bottom_right({trees[474], lumberyards[474]}), .init(2'b00), .state({trees[423], lumberyards[423]}));
acre acre_8_24 (.clk(clk), .en(en), .top_left({trees[373], lumberyards[373]}), .top({trees[374], lumberyards[374]}), .top_right({trees[375], lumberyards[375]}), .left({trees[423], lumberyards[423]}), .right({trees[425], lumberyards[425]}), .bottom_left({trees[473], lumberyards[473]}), .bottom({trees[474], lumberyards[474]}), .bottom_right({trees[475], lumberyards[475]}), .init(2'b10), .state({trees[424], lumberyards[424]}));
acre acre_8_25 (.clk(clk), .en(en), .top_left({trees[374], lumberyards[374]}), .top({trees[375], lumberyards[375]}), .top_right({trees[376], lumberyards[376]}), .left({trees[424], lumberyards[424]}), .right({trees[426], lumberyards[426]}), .bottom_left({trees[474], lumberyards[474]}), .bottom({trees[475], lumberyards[475]}), .bottom_right({trees[476], lumberyards[476]}), .init(2'b00), .state({trees[425], lumberyards[425]}));
acre acre_8_26 (.clk(clk), .en(en), .top_left({trees[375], lumberyards[375]}), .top({trees[376], lumberyards[376]}), .top_right({trees[377], lumberyards[377]}), .left({trees[425], lumberyards[425]}), .right({trees[427], lumberyards[427]}), .bottom_left({trees[475], lumberyards[475]}), .bottom({trees[476], lumberyards[476]}), .bottom_right({trees[477], lumberyards[477]}), .init(2'b00), .state({trees[426], lumberyards[426]}));
acre acre_8_27 (.clk(clk), .en(en), .top_left({trees[376], lumberyards[376]}), .top({trees[377], lumberyards[377]}), .top_right({trees[378], lumberyards[378]}), .left({trees[426], lumberyards[426]}), .right({trees[428], lumberyards[428]}), .bottom_left({trees[476], lumberyards[476]}), .bottom({trees[477], lumberyards[477]}), .bottom_right({trees[478], lumberyards[478]}), .init(2'b00), .state({trees[427], lumberyards[427]}));
acre acre_8_28 (.clk(clk), .en(en), .top_left({trees[377], lumberyards[377]}), .top({trees[378], lumberyards[378]}), .top_right({trees[379], lumberyards[379]}), .left({trees[427], lumberyards[427]}), .right({trees[429], lumberyards[429]}), .bottom_left({trees[477], lumberyards[477]}), .bottom({trees[478], lumberyards[478]}), .bottom_right({trees[479], lumberyards[479]}), .init(2'b00), .state({trees[428], lumberyards[428]}));
acre acre_8_29 (.clk(clk), .en(en), .top_left({trees[378], lumberyards[378]}), .top({trees[379], lumberyards[379]}), .top_right({trees[380], lumberyards[380]}), .left({trees[428], lumberyards[428]}), .right({trees[430], lumberyards[430]}), .bottom_left({trees[478], lumberyards[478]}), .bottom({trees[479], lumberyards[479]}), .bottom_right({trees[480], lumberyards[480]}), .init(2'b00), .state({trees[429], lumberyards[429]}));
acre acre_8_30 (.clk(clk), .en(en), .top_left({trees[379], lumberyards[379]}), .top({trees[380], lumberyards[380]}), .top_right({trees[381], lumberyards[381]}), .left({trees[429], lumberyards[429]}), .right({trees[431], lumberyards[431]}), .bottom_left({trees[479], lumberyards[479]}), .bottom({trees[480], lumberyards[480]}), .bottom_right({trees[481], lumberyards[481]}), .init(2'b00), .state({trees[430], lumberyards[430]}));
acre acre_8_31 (.clk(clk), .en(en), .top_left({trees[380], lumberyards[380]}), .top({trees[381], lumberyards[381]}), .top_right({trees[382], lumberyards[382]}), .left({trees[430], lumberyards[430]}), .right({trees[432], lumberyards[432]}), .bottom_left({trees[480], lumberyards[480]}), .bottom({trees[481], lumberyards[481]}), .bottom_right({trees[482], lumberyards[482]}), .init(2'b00), .state({trees[431], lumberyards[431]}));
acre acre_8_32 (.clk(clk), .en(en), .top_left({trees[381], lumberyards[381]}), .top({trees[382], lumberyards[382]}), .top_right({trees[383], lumberyards[383]}), .left({trees[431], lumberyards[431]}), .right({trees[433], lumberyards[433]}), .bottom_left({trees[481], lumberyards[481]}), .bottom({trees[482], lumberyards[482]}), .bottom_right({trees[483], lumberyards[483]}), .init(2'b10), .state({trees[432], lumberyards[432]}));
acre acre_8_33 (.clk(clk), .en(en), .top_left({trees[382], lumberyards[382]}), .top({trees[383], lumberyards[383]}), .top_right({trees[384], lumberyards[384]}), .left({trees[432], lumberyards[432]}), .right({trees[434], lumberyards[434]}), .bottom_left({trees[482], lumberyards[482]}), .bottom({trees[483], lumberyards[483]}), .bottom_right({trees[484], lumberyards[484]}), .init(2'b00), .state({trees[433], lumberyards[433]}));
acre acre_8_34 (.clk(clk), .en(en), .top_left({trees[383], lumberyards[383]}), .top({trees[384], lumberyards[384]}), .top_right({trees[385], lumberyards[385]}), .left({trees[433], lumberyards[433]}), .right({trees[435], lumberyards[435]}), .bottom_left({trees[483], lumberyards[483]}), .bottom({trees[484], lumberyards[484]}), .bottom_right({trees[485], lumberyards[485]}), .init(2'b01), .state({trees[434], lumberyards[434]}));
acre acre_8_35 (.clk(clk), .en(en), .top_left({trees[384], lumberyards[384]}), .top({trees[385], lumberyards[385]}), .top_right({trees[386], lumberyards[386]}), .left({trees[434], lumberyards[434]}), .right({trees[436], lumberyards[436]}), .bottom_left({trees[484], lumberyards[484]}), .bottom({trees[485], lumberyards[485]}), .bottom_right({trees[486], lumberyards[486]}), .init(2'b00), .state({trees[435], lumberyards[435]}));
acre acre_8_36 (.clk(clk), .en(en), .top_left({trees[385], lumberyards[385]}), .top({trees[386], lumberyards[386]}), .top_right({trees[387], lumberyards[387]}), .left({trees[435], lumberyards[435]}), .right({trees[437], lumberyards[437]}), .bottom_left({trees[485], lumberyards[485]}), .bottom({trees[486], lumberyards[486]}), .bottom_right({trees[487], lumberyards[487]}), .init(2'b00), .state({trees[436], lumberyards[436]}));
acre acre_8_37 (.clk(clk), .en(en), .top_left({trees[386], lumberyards[386]}), .top({trees[387], lumberyards[387]}), .top_right({trees[388], lumberyards[388]}), .left({trees[436], lumberyards[436]}), .right({trees[438], lumberyards[438]}), .bottom_left({trees[486], lumberyards[486]}), .bottom({trees[487], lumberyards[487]}), .bottom_right({trees[488], lumberyards[488]}), .init(2'b10), .state({trees[437], lumberyards[437]}));
acre acre_8_38 (.clk(clk), .en(en), .top_left({trees[387], lumberyards[387]}), .top({trees[388], lumberyards[388]}), .top_right({trees[389], lumberyards[389]}), .left({trees[437], lumberyards[437]}), .right({trees[439], lumberyards[439]}), .bottom_left({trees[487], lumberyards[487]}), .bottom({trees[488], lumberyards[488]}), .bottom_right({trees[489], lumberyards[489]}), .init(2'b00), .state({trees[438], lumberyards[438]}));
acre acre_8_39 (.clk(clk), .en(en), .top_left({trees[388], lumberyards[388]}), .top({trees[389], lumberyards[389]}), .top_right({trees[390], lumberyards[390]}), .left({trees[438], lumberyards[438]}), .right({trees[440], lumberyards[440]}), .bottom_left({trees[488], lumberyards[488]}), .bottom({trees[489], lumberyards[489]}), .bottom_right({trees[490], lumberyards[490]}), .init(2'b00), .state({trees[439], lumberyards[439]}));
acre acre_8_40 (.clk(clk), .en(en), .top_left({trees[389], lumberyards[389]}), .top({trees[390], lumberyards[390]}), .top_right({trees[391], lumberyards[391]}), .left({trees[439], lumberyards[439]}), .right({trees[441], lumberyards[441]}), .bottom_left({trees[489], lumberyards[489]}), .bottom({trees[490], lumberyards[490]}), .bottom_right({trees[491], lumberyards[491]}), .init(2'b00), .state({trees[440], lumberyards[440]}));
acre acre_8_41 (.clk(clk), .en(en), .top_left({trees[390], lumberyards[390]}), .top({trees[391], lumberyards[391]}), .top_right({trees[392], lumberyards[392]}), .left({trees[440], lumberyards[440]}), .right({trees[442], lumberyards[442]}), .bottom_left({trees[490], lumberyards[490]}), .bottom({trees[491], lumberyards[491]}), .bottom_right({trees[492], lumberyards[492]}), .init(2'b00), .state({trees[441], lumberyards[441]}));
acre acre_8_42 (.clk(clk), .en(en), .top_left({trees[391], lumberyards[391]}), .top({trees[392], lumberyards[392]}), .top_right({trees[393], lumberyards[393]}), .left({trees[441], lumberyards[441]}), .right({trees[443], lumberyards[443]}), .bottom_left({trees[491], lumberyards[491]}), .bottom({trees[492], lumberyards[492]}), .bottom_right({trees[493], lumberyards[493]}), .init(2'b00), .state({trees[442], lumberyards[442]}));
acre acre_8_43 (.clk(clk), .en(en), .top_left({trees[392], lumberyards[392]}), .top({trees[393], lumberyards[393]}), .top_right({trees[394], lumberyards[394]}), .left({trees[442], lumberyards[442]}), .right({trees[444], lumberyards[444]}), .bottom_left({trees[492], lumberyards[492]}), .bottom({trees[493], lumberyards[493]}), .bottom_right({trees[494], lumberyards[494]}), .init(2'b00), .state({trees[443], lumberyards[443]}));
acre acre_8_44 (.clk(clk), .en(en), .top_left({trees[393], lumberyards[393]}), .top({trees[394], lumberyards[394]}), .top_right({trees[395], lumberyards[395]}), .left({trees[443], lumberyards[443]}), .right({trees[445], lumberyards[445]}), .bottom_left({trees[493], lumberyards[493]}), .bottom({trees[494], lumberyards[494]}), .bottom_right({trees[495], lumberyards[495]}), .init(2'b00), .state({trees[444], lumberyards[444]}));
acre acre_8_45 (.clk(clk), .en(en), .top_left({trees[394], lumberyards[394]}), .top({trees[395], lumberyards[395]}), .top_right({trees[396], lumberyards[396]}), .left({trees[444], lumberyards[444]}), .right({trees[446], lumberyards[446]}), .bottom_left({trees[494], lumberyards[494]}), .bottom({trees[495], lumberyards[495]}), .bottom_right({trees[496], lumberyards[496]}), .init(2'b01), .state({trees[445], lumberyards[445]}));
acre acre_8_46 (.clk(clk), .en(en), .top_left({trees[395], lumberyards[395]}), .top({trees[396], lumberyards[396]}), .top_right({trees[397], lumberyards[397]}), .left({trees[445], lumberyards[445]}), .right({trees[447], lumberyards[447]}), .bottom_left({trees[495], lumberyards[495]}), .bottom({trees[496], lumberyards[496]}), .bottom_right({trees[497], lumberyards[497]}), .init(2'b10), .state({trees[446], lumberyards[446]}));
acre acre_8_47 (.clk(clk), .en(en), .top_left({trees[396], lumberyards[396]}), .top({trees[397], lumberyards[397]}), .top_right({trees[398], lumberyards[398]}), .left({trees[446], lumberyards[446]}), .right({trees[448], lumberyards[448]}), .bottom_left({trees[496], lumberyards[496]}), .bottom({trees[497], lumberyards[497]}), .bottom_right({trees[498], lumberyards[498]}), .init(2'b00), .state({trees[447], lumberyards[447]}));
acre acre_8_48 (.clk(clk), .en(en), .top_left({trees[397], lumberyards[397]}), .top({trees[398], lumberyards[398]}), .top_right({trees[399], lumberyards[399]}), .left({trees[447], lumberyards[447]}), .right({trees[449], lumberyards[449]}), .bottom_left({trees[497], lumberyards[497]}), .bottom({trees[498], lumberyards[498]}), .bottom_right({trees[499], lumberyards[499]}), .init(2'b10), .state({trees[448], lumberyards[448]}));
acre acre_8_49 (.clk(clk), .en(en), .top_left({trees[398], lumberyards[398]}), .top({trees[399], lumberyards[399]}), .top_right(2'b0), .left({trees[448], lumberyards[448]}), .right(2'b0), .bottom_left({trees[498], lumberyards[498]}), .bottom({trees[499], lumberyards[499]}), .bottom_right(2'b0), .init(2'b00), .state({trees[449], lumberyards[449]}));
acre acre_9_0 (.clk(clk), .en(en), .top_left(2'b0), .top({trees[400], lumberyards[400]}), .top_right({trees[401], lumberyards[401]}), .left(2'b0), .right({trees[451], lumberyards[451]}), .bottom_left(2'b0), .bottom({trees[500], lumberyards[500]}), .bottom_right({trees[501], lumberyards[501]}), .init(2'b00), .state({trees[450], lumberyards[450]}));
acre acre_9_1 (.clk(clk), .en(en), .top_left({trees[400], lumberyards[400]}), .top({trees[401], lumberyards[401]}), .top_right({trees[402], lumberyards[402]}), .left({trees[450], lumberyards[450]}), .right({trees[452], lumberyards[452]}), .bottom_left({trees[500], lumberyards[500]}), .bottom({trees[501], lumberyards[501]}), .bottom_right({trees[502], lumberyards[502]}), .init(2'b00), .state({trees[451], lumberyards[451]}));
acre acre_9_2 (.clk(clk), .en(en), .top_left({trees[401], lumberyards[401]}), .top({trees[402], lumberyards[402]}), .top_right({trees[403], lumberyards[403]}), .left({trees[451], lumberyards[451]}), .right({trees[453], lumberyards[453]}), .bottom_left({trees[501], lumberyards[501]}), .bottom({trees[502], lumberyards[502]}), .bottom_right({trees[503], lumberyards[503]}), .init(2'b00), .state({trees[452], lumberyards[452]}));
acre acre_9_3 (.clk(clk), .en(en), .top_left({trees[402], lumberyards[402]}), .top({trees[403], lumberyards[403]}), .top_right({trees[404], lumberyards[404]}), .left({trees[452], lumberyards[452]}), .right({trees[454], lumberyards[454]}), .bottom_left({trees[502], lumberyards[502]}), .bottom({trees[503], lumberyards[503]}), .bottom_right({trees[504], lumberyards[504]}), .init(2'b10), .state({trees[453], lumberyards[453]}));
acre acre_9_4 (.clk(clk), .en(en), .top_left({trees[403], lumberyards[403]}), .top({trees[404], lumberyards[404]}), .top_right({trees[405], lumberyards[405]}), .left({trees[453], lumberyards[453]}), .right({trees[455], lumberyards[455]}), .bottom_left({trees[503], lumberyards[503]}), .bottom({trees[504], lumberyards[504]}), .bottom_right({trees[505], lumberyards[505]}), .init(2'b00), .state({trees[454], lumberyards[454]}));
acre acre_9_5 (.clk(clk), .en(en), .top_left({trees[404], lumberyards[404]}), .top({trees[405], lumberyards[405]}), .top_right({trees[406], lumberyards[406]}), .left({trees[454], lumberyards[454]}), .right({trees[456], lumberyards[456]}), .bottom_left({trees[504], lumberyards[504]}), .bottom({trees[505], lumberyards[505]}), .bottom_right({trees[506], lumberyards[506]}), .init(2'b10), .state({trees[455], lumberyards[455]}));
acre acre_9_6 (.clk(clk), .en(en), .top_left({trees[405], lumberyards[405]}), .top({trees[406], lumberyards[406]}), .top_right({trees[407], lumberyards[407]}), .left({trees[455], lumberyards[455]}), .right({trees[457], lumberyards[457]}), .bottom_left({trees[505], lumberyards[505]}), .bottom({trees[506], lumberyards[506]}), .bottom_right({trees[507], lumberyards[507]}), .init(2'b01), .state({trees[456], lumberyards[456]}));
acre acre_9_7 (.clk(clk), .en(en), .top_left({trees[406], lumberyards[406]}), .top({trees[407], lumberyards[407]}), .top_right({trees[408], lumberyards[408]}), .left({trees[456], lumberyards[456]}), .right({trees[458], lumberyards[458]}), .bottom_left({trees[506], lumberyards[506]}), .bottom({trees[507], lumberyards[507]}), .bottom_right({trees[508], lumberyards[508]}), .init(2'b00), .state({trees[457], lumberyards[457]}));
acre acre_9_8 (.clk(clk), .en(en), .top_left({trees[407], lumberyards[407]}), .top({trees[408], lumberyards[408]}), .top_right({trees[409], lumberyards[409]}), .left({trees[457], lumberyards[457]}), .right({trees[459], lumberyards[459]}), .bottom_left({trees[507], lumberyards[507]}), .bottom({trees[508], lumberyards[508]}), .bottom_right({trees[509], lumberyards[509]}), .init(2'b00), .state({trees[458], lumberyards[458]}));
acre acre_9_9 (.clk(clk), .en(en), .top_left({trees[408], lumberyards[408]}), .top({trees[409], lumberyards[409]}), .top_right({trees[410], lumberyards[410]}), .left({trees[458], lumberyards[458]}), .right({trees[460], lumberyards[460]}), .bottom_left({trees[508], lumberyards[508]}), .bottom({trees[509], lumberyards[509]}), .bottom_right({trees[510], lumberyards[510]}), .init(2'b10), .state({trees[459], lumberyards[459]}));
acre acre_9_10 (.clk(clk), .en(en), .top_left({trees[409], lumberyards[409]}), .top({trees[410], lumberyards[410]}), .top_right({trees[411], lumberyards[411]}), .left({trees[459], lumberyards[459]}), .right({trees[461], lumberyards[461]}), .bottom_left({trees[509], lumberyards[509]}), .bottom({trees[510], lumberyards[510]}), .bottom_right({trees[511], lumberyards[511]}), .init(2'b00), .state({trees[460], lumberyards[460]}));
acre acre_9_11 (.clk(clk), .en(en), .top_left({trees[410], lumberyards[410]}), .top({trees[411], lumberyards[411]}), .top_right({trees[412], lumberyards[412]}), .left({trees[460], lumberyards[460]}), .right({trees[462], lumberyards[462]}), .bottom_left({trees[510], lumberyards[510]}), .bottom({trees[511], lumberyards[511]}), .bottom_right({trees[512], lumberyards[512]}), .init(2'b00), .state({trees[461], lumberyards[461]}));
acre acre_9_12 (.clk(clk), .en(en), .top_left({trees[411], lumberyards[411]}), .top({trees[412], lumberyards[412]}), .top_right({trees[413], lumberyards[413]}), .left({trees[461], lumberyards[461]}), .right({trees[463], lumberyards[463]}), .bottom_left({trees[511], lumberyards[511]}), .bottom({trees[512], lumberyards[512]}), .bottom_right({trees[513], lumberyards[513]}), .init(2'b00), .state({trees[462], lumberyards[462]}));
acre acre_9_13 (.clk(clk), .en(en), .top_left({trees[412], lumberyards[412]}), .top({trees[413], lumberyards[413]}), .top_right({trees[414], lumberyards[414]}), .left({trees[462], lumberyards[462]}), .right({trees[464], lumberyards[464]}), .bottom_left({trees[512], lumberyards[512]}), .bottom({trees[513], lumberyards[513]}), .bottom_right({trees[514], lumberyards[514]}), .init(2'b00), .state({trees[463], lumberyards[463]}));
acre acre_9_14 (.clk(clk), .en(en), .top_left({trees[413], lumberyards[413]}), .top({trees[414], lumberyards[414]}), .top_right({trees[415], lumberyards[415]}), .left({trees[463], lumberyards[463]}), .right({trees[465], lumberyards[465]}), .bottom_left({trees[513], lumberyards[513]}), .bottom({trees[514], lumberyards[514]}), .bottom_right({trees[515], lumberyards[515]}), .init(2'b10), .state({trees[464], lumberyards[464]}));
acre acre_9_15 (.clk(clk), .en(en), .top_left({trees[414], lumberyards[414]}), .top({trees[415], lumberyards[415]}), .top_right({trees[416], lumberyards[416]}), .left({trees[464], lumberyards[464]}), .right({trees[466], lumberyards[466]}), .bottom_left({trees[514], lumberyards[514]}), .bottom({trees[515], lumberyards[515]}), .bottom_right({trees[516], lumberyards[516]}), .init(2'b00), .state({trees[465], lumberyards[465]}));
acre acre_9_16 (.clk(clk), .en(en), .top_left({trees[415], lumberyards[415]}), .top({trees[416], lumberyards[416]}), .top_right({trees[417], lumberyards[417]}), .left({trees[465], lumberyards[465]}), .right({trees[467], lumberyards[467]}), .bottom_left({trees[515], lumberyards[515]}), .bottom({trees[516], lumberyards[516]}), .bottom_right({trees[517], lumberyards[517]}), .init(2'b00), .state({trees[466], lumberyards[466]}));
acre acre_9_17 (.clk(clk), .en(en), .top_left({trees[416], lumberyards[416]}), .top({trees[417], lumberyards[417]}), .top_right({trees[418], lumberyards[418]}), .left({trees[466], lumberyards[466]}), .right({trees[468], lumberyards[468]}), .bottom_left({trees[516], lumberyards[516]}), .bottom({trees[517], lumberyards[517]}), .bottom_right({trees[518], lumberyards[518]}), .init(2'b00), .state({trees[467], lumberyards[467]}));
acre acre_9_18 (.clk(clk), .en(en), .top_left({trees[417], lumberyards[417]}), .top({trees[418], lumberyards[418]}), .top_right({trees[419], lumberyards[419]}), .left({trees[467], lumberyards[467]}), .right({trees[469], lumberyards[469]}), .bottom_left({trees[517], lumberyards[517]}), .bottom({trees[518], lumberyards[518]}), .bottom_right({trees[519], lumberyards[519]}), .init(2'b00), .state({trees[468], lumberyards[468]}));
acre acre_9_19 (.clk(clk), .en(en), .top_left({trees[418], lumberyards[418]}), .top({trees[419], lumberyards[419]}), .top_right({trees[420], lumberyards[420]}), .left({trees[468], lumberyards[468]}), .right({trees[470], lumberyards[470]}), .bottom_left({trees[518], lumberyards[518]}), .bottom({trees[519], lumberyards[519]}), .bottom_right({trees[520], lumberyards[520]}), .init(2'b01), .state({trees[469], lumberyards[469]}));
acre acre_9_20 (.clk(clk), .en(en), .top_left({trees[419], lumberyards[419]}), .top({trees[420], lumberyards[420]}), .top_right({trees[421], lumberyards[421]}), .left({trees[469], lumberyards[469]}), .right({trees[471], lumberyards[471]}), .bottom_left({trees[519], lumberyards[519]}), .bottom({trees[520], lumberyards[520]}), .bottom_right({trees[521], lumberyards[521]}), .init(2'b00), .state({trees[470], lumberyards[470]}));
acre acre_9_21 (.clk(clk), .en(en), .top_left({trees[420], lumberyards[420]}), .top({trees[421], lumberyards[421]}), .top_right({trees[422], lumberyards[422]}), .left({trees[470], lumberyards[470]}), .right({trees[472], lumberyards[472]}), .bottom_left({trees[520], lumberyards[520]}), .bottom({trees[521], lumberyards[521]}), .bottom_right({trees[522], lumberyards[522]}), .init(2'b00), .state({trees[471], lumberyards[471]}));
acre acre_9_22 (.clk(clk), .en(en), .top_left({trees[421], lumberyards[421]}), .top({trees[422], lumberyards[422]}), .top_right({trees[423], lumberyards[423]}), .left({trees[471], lumberyards[471]}), .right({trees[473], lumberyards[473]}), .bottom_left({trees[521], lumberyards[521]}), .bottom({trees[522], lumberyards[522]}), .bottom_right({trees[523], lumberyards[523]}), .init(2'b10), .state({trees[472], lumberyards[472]}));
acre acre_9_23 (.clk(clk), .en(en), .top_left({trees[422], lumberyards[422]}), .top({trees[423], lumberyards[423]}), .top_right({trees[424], lumberyards[424]}), .left({trees[472], lumberyards[472]}), .right({trees[474], lumberyards[474]}), .bottom_left({trees[522], lumberyards[522]}), .bottom({trees[523], lumberyards[523]}), .bottom_right({trees[524], lumberyards[524]}), .init(2'b10), .state({trees[473], lumberyards[473]}));
acre acre_9_24 (.clk(clk), .en(en), .top_left({trees[423], lumberyards[423]}), .top({trees[424], lumberyards[424]}), .top_right({trees[425], lumberyards[425]}), .left({trees[473], lumberyards[473]}), .right({trees[475], lumberyards[475]}), .bottom_left({trees[523], lumberyards[523]}), .bottom({trees[524], lumberyards[524]}), .bottom_right({trees[525], lumberyards[525]}), .init(2'b01), .state({trees[474], lumberyards[474]}));
acre acre_9_25 (.clk(clk), .en(en), .top_left({trees[424], lumberyards[424]}), .top({trees[425], lumberyards[425]}), .top_right({trees[426], lumberyards[426]}), .left({trees[474], lumberyards[474]}), .right({trees[476], lumberyards[476]}), .bottom_left({trees[524], lumberyards[524]}), .bottom({trees[525], lumberyards[525]}), .bottom_right({trees[526], lumberyards[526]}), .init(2'b00), .state({trees[475], lumberyards[475]}));
acre acre_9_26 (.clk(clk), .en(en), .top_left({trees[425], lumberyards[425]}), .top({trees[426], lumberyards[426]}), .top_right({trees[427], lumberyards[427]}), .left({trees[475], lumberyards[475]}), .right({trees[477], lumberyards[477]}), .bottom_left({trees[525], lumberyards[525]}), .bottom({trees[526], lumberyards[526]}), .bottom_right({trees[527], lumberyards[527]}), .init(2'b10), .state({trees[476], lumberyards[476]}));
acre acre_9_27 (.clk(clk), .en(en), .top_left({trees[426], lumberyards[426]}), .top({trees[427], lumberyards[427]}), .top_right({trees[428], lumberyards[428]}), .left({trees[476], lumberyards[476]}), .right({trees[478], lumberyards[478]}), .bottom_left({trees[526], lumberyards[526]}), .bottom({trees[527], lumberyards[527]}), .bottom_right({trees[528], lumberyards[528]}), .init(2'b00), .state({trees[477], lumberyards[477]}));
acre acre_9_28 (.clk(clk), .en(en), .top_left({trees[427], lumberyards[427]}), .top({trees[428], lumberyards[428]}), .top_right({trees[429], lumberyards[429]}), .left({trees[477], lumberyards[477]}), .right({trees[479], lumberyards[479]}), .bottom_left({trees[527], lumberyards[527]}), .bottom({trees[528], lumberyards[528]}), .bottom_right({trees[529], lumberyards[529]}), .init(2'b01), .state({trees[478], lumberyards[478]}));
acre acre_9_29 (.clk(clk), .en(en), .top_left({trees[428], lumberyards[428]}), .top({trees[429], lumberyards[429]}), .top_right({trees[430], lumberyards[430]}), .left({trees[478], lumberyards[478]}), .right({trees[480], lumberyards[480]}), .bottom_left({trees[528], lumberyards[528]}), .bottom({trees[529], lumberyards[529]}), .bottom_right({trees[530], lumberyards[530]}), .init(2'b00), .state({trees[479], lumberyards[479]}));
acre acre_9_30 (.clk(clk), .en(en), .top_left({trees[429], lumberyards[429]}), .top({trees[430], lumberyards[430]}), .top_right({trees[431], lumberyards[431]}), .left({trees[479], lumberyards[479]}), .right({trees[481], lumberyards[481]}), .bottom_left({trees[529], lumberyards[529]}), .bottom({trees[530], lumberyards[530]}), .bottom_right({trees[531], lumberyards[531]}), .init(2'b00), .state({trees[480], lumberyards[480]}));
acre acre_9_31 (.clk(clk), .en(en), .top_left({trees[430], lumberyards[430]}), .top({trees[431], lumberyards[431]}), .top_right({trees[432], lumberyards[432]}), .left({trees[480], lumberyards[480]}), .right({trees[482], lumberyards[482]}), .bottom_left({trees[530], lumberyards[530]}), .bottom({trees[531], lumberyards[531]}), .bottom_right({trees[532], lumberyards[532]}), .init(2'b10), .state({trees[481], lumberyards[481]}));
acre acre_9_32 (.clk(clk), .en(en), .top_left({trees[431], lumberyards[431]}), .top({trees[432], lumberyards[432]}), .top_right({trees[433], lumberyards[433]}), .left({trees[481], lumberyards[481]}), .right({trees[483], lumberyards[483]}), .bottom_left({trees[531], lumberyards[531]}), .bottom({trees[532], lumberyards[532]}), .bottom_right({trees[533], lumberyards[533]}), .init(2'b00), .state({trees[482], lumberyards[482]}));
acre acre_9_33 (.clk(clk), .en(en), .top_left({trees[432], lumberyards[432]}), .top({trees[433], lumberyards[433]}), .top_right({trees[434], lumberyards[434]}), .left({trees[482], lumberyards[482]}), .right({trees[484], lumberyards[484]}), .bottom_left({trees[532], lumberyards[532]}), .bottom({trees[533], lumberyards[533]}), .bottom_right({trees[534], lumberyards[534]}), .init(2'b00), .state({trees[483], lumberyards[483]}));
acre acre_9_34 (.clk(clk), .en(en), .top_left({trees[433], lumberyards[433]}), .top({trees[434], lumberyards[434]}), .top_right({trees[435], lumberyards[435]}), .left({trees[483], lumberyards[483]}), .right({trees[485], lumberyards[485]}), .bottom_left({trees[533], lumberyards[533]}), .bottom({trees[534], lumberyards[534]}), .bottom_right({trees[535], lumberyards[535]}), .init(2'b00), .state({trees[484], lumberyards[484]}));
acre acre_9_35 (.clk(clk), .en(en), .top_left({trees[434], lumberyards[434]}), .top({trees[435], lumberyards[435]}), .top_right({trees[436], lumberyards[436]}), .left({trees[484], lumberyards[484]}), .right({trees[486], lumberyards[486]}), .bottom_left({trees[534], lumberyards[534]}), .bottom({trees[535], lumberyards[535]}), .bottom_right({trees[536], lumberyards[536]}), .init(2'b00), .state({trees[485], lumberyards[485]}));
acre acre_9_36 (.clk(clk), .en(en), .top_left({trees[435], lumberyards[435]}), .top({trees[436], lumberyards[436]}), .top_right({trees[437], lumberyards[437]}), .left({trees[485], lumberyards[485]}), .right({trees[487], lumberyards[487]}), .bottom_left({trees[535], lumberyards[535]}), .bottom({trees[536], lumberyards[536]}), .bottom_right({trees[537], lumberyards[537]}), .init(2'b00), .state({trees[486], lumberyards[486]}));
acre acre_9_37 (.clk(clk), .en(en), .top_left({trees[436], lumberyards[436]}), .top({trees[437], lumberyards[437]}), .top_right({trees[438], lumberyards[438]}), .left({trees[486], lumberyards[486]}), .right({trees[488], lumberyards[488]}), .bottom_left({trees[536], lumberyards[536]}), .bottom({trees[537], lumberyards[537]}), .bottom_right({trees[538], lumberyards[538]}), .init(2'b10), .state({trees[487], lumberyards[487]}));
acre acre_9_38 (.clk(clk), .en(en), .top_left({trees[437], lumberyards[437]}), .top({trees[438], lumberyards[438]}), .top_right({trees[439], lumberyards[439]}), .left({trees[487], lumberyards[487]}), .right({trees[489], lumberyards[489]}), .bottom_left({trees[537], lumberyards[537]}), .bottom({trees[538], lumberyards[538]}), .bottom_right({trees[539], lumberyards[539]}), .init(2'b00), .state({trees[488], lumberyards[488]}));
acre acre_9_39 (.clk(clk), .en(en), .top_left({trees[438], lumberyards[438]}), .top({trees[439], lumberyards[439]}), .top_right({trees[440], lumberyards[440]}), .left({trees[488], lumberyards[488]}), .right({trees[490], lumberyards[490]}), .bottom_left({trees[538], lumberyards[538]}), .bottom({trees[539], lumberyards[539]}), .bottom_right({trees[540], lumberyards[540]}), .init(2'b00), .state({trees[489], lumberyards[489]}));
acre acre_9_40 (.clk(clk), .en(en), .top_left({trees[439], lumberyards[439]}), .top({trees[440], lumberyards[440]}), .top_right({trees[441], lumberyards[441]}), .left({trees[489], lumberyards[489]}), .right({trees[491], lumberyards[491]}), .bottom_left({trees[539], lumberyards[539]}), .bottom({trees[540], lumberyards[540]}), .bottom_right({trees[541], lumberyards[541]}), .init(2'b01), .state({trees[490], lumberyards[490]}));
acre acre_9_41 (.clk(clk), .en(en), .top_left({trees[440], lumberyards[440]}), .top({trees[441], lumberyards[441]}), .top_right({trees[442], lumberyards[442]}), .left({trees[490], lumberyards[490]}), .right({trees[492], lumberyards[492]}), .bottom_left({trees[540], lumberyards[540]}), .bottom({trees[541], lumberyards[541]}), .bottom_right({trees[542], lumberyards[542]}), .init(2'b00), .state({trees[491], lumberyards[491]}));
acre acre_9_42 (.clk(clk), .en(en), .top_left({trees[441], lumberyards[441]}), .top({trees[442], lumberyards[442]}), .top_right({trees[443], lumberyards[443]}), .left({trees[491], lumberyards[491]}), .right({trees[493], lumberyards[493]}), .bottom_left({trees[541], lumberyards[541]}), .bottom({trees[542], lumberyards[542]}), .bottom_right({trees[543], lumberyards[543]}), .init(2'b00), .state({trees[492], lumberyards[492]}));
acre acre_9_43 (.clk(clk), .en(en), .top_left({trees[442], lumberyards[442]}), .top({trees[443], lumberyards[443]}), .top_right({trees[444], lumberyards[444]}), .left({trees[492], lumberyards[492]}), .right({trees[494], lumberyards[494]}), .bottom_left({trees[542], lumberyards[542]}), .bottom({trees[543], lumberyards[543]}), .bottom_right({trees[544], lumberyards[544]}), .init(2'b00), .state({trees[493], lumberyards[493]}));
acre acre_9_44 (.clk(clk), .en(en), .top_left({trees[443], lumberyards[443]}), .top({trees[444], lumberyards[444]}), .top_right({trees[445], lumberyards[445]}), .left({trees[493], lumberyards[493]}), .right({trees[495], lumberyards[495]}), .bottom_left({trees[543], lumberyards[543]}), .bottom({trees[544], lumberyards[544]}), .bottom_right({trees[545], lumberyards[545]}), .init(2'b00), .state({trees[494], lumberyards[494]}));
acre acre_9_45 (.clk(clk), .en(en), .top_left({trees[444], lumberyards[444]}), .top({trees[445], lumberyards[445]}), .top_right({trees[446], lumberyards[446]}), .left({trees[494], lumberyards[494]}), .right({trees[496], lumberyards[496]}), .bottom_left({trees[544], lumberyards[544]}), .bottom({trees[545], lumberyards[545]}), .bottom_right({trees[546], lumberyards[546]}), .init(2'b00), .state({trees[495], lumberyards[495]}));
acre acre_9_46 (.clk(clk), .en(en), .top_left({trees[445], lumberyards[445]}), .top({trees[446], lumberyards[446]}), .top_right({trees[447], lumberyards[447]}), .left({trees[495], lumberyards[495]}), .right({trees[497], lumberyards[497]}), .bottom_left({trees[545], lumberyards[545]}), .bottom({trees[546], lumberyards[546]}), .bottom_right({trees[547], lumberyards[547]}), .init(2'b01), .state({trees[496], lumberyards[496]}));
acre acre_9_47 (.clk(clk), .en(en), .top_left({trees[446], lumberyards[446]}), .top({trees[447], lumberyards[447]}), .top_right({trees[448], lumberyards[448]}), .left({trees[496], lumberyards[496]}), .right({trees[498], lumberyards[498]}), .bottom_left({trees[546], lumberyards[546]}), .bottom({trees[547], lumberyards[547]}), .bottom_right({trees[548], lumberyards[548]}), .init(2'b00), .state({trees[497], lumberyards[497]}));
acre acre_9_48 (.clk(clk), .en(en), .top_left({trees[447], lumberyards[447]}), .top({trees[448], lumberyards[448]}), .top_right({trees[449], lumberyards[449]}), .left({trees[497], lumberyards[497]}), .right({trees[499], lumberyards[499]}), .bottom_left({trees[547], lumberyards[547]}), .bottom({trees[548], lumberyards[548]}), .bottom_right({trees[549], lumberyards[549]}), .init(2'b00), .state({trees[498], lumberyards[498]}));
acre acre_9_49 (.clk(clk), .en(en), .top_left({trees[448], lumberyards[448]}), .top({trees[449], lumberyards[449]}), .top_right(2'b0), .left({trees[498], lumberyards[498]}), .right(2'b0), .bottom_left({trees[548], lumberyards[548]}), .bottom({trees[549], lumberyards[549]}), .bottom_right(2'b0), .init(2'b00), .state({trees[499], lumberyards[499]}));
acre acre_10_0 (.clk(clk), .en(en), .top_left(2'b0), .top({trees[450], lumberyards[450]}), .top_right({trees[451], lumberyards[451]}), .left(2'b0), .right({trees[501], lumberyards[501]}), .bottom_left(2'b0), .bottom({trees[550], lumberyards[550]}), .bottom_right({trees[551], lumberyards[551]}), .init(2'b00), .state({trees[500], lumberyards[500]}));
acre acre_10_1 (.clk(clk), .en(en), .top_left({trees[450], lumberyards[450]}), .top({trees[451], lumberyards[451]}), .top_right({trees[452], lumberyards[452]}), .left({trees[500], lumberyards[500]}), .right({trees[502], lumberyards[502]}), .bottom_left({trees[550], lumberyards[550]}), .bottom({trees[551], lumberyards[551]}), .bottom_right({trees[552], lumberyards[552]}), .init(2'b10), .state({trees[501], lumberyards[501]}));
acre acre_10_2 (.clk(clk), .en(en), .top_left({trees[451], lumberyards[451]}), .top({trees[452], lumberyards[452]}), .top_right({trees[453], lumberyards[453]}), .left({trees[501], lumberyards[501]}), .right({trees[503], lumberyards[503]}), .bottom_left({trees[551], lumberyards[551]}), .bottom({trees[552], lumberyards[552]}), .bottom_right({trees[553], lumberyards[553]}), .init(2'b00), .state({trees[502], lumberyards[502]}));
acre acre_10_3 (.clk(clk), .en(en), .top_left({trees[452], lumberyards[452]}), .top({trees[453], lumberyards[453]}), .top_right({trees[454], lumberyards[454]}), .left({trees[502], lumberyards[502]}), .right({trees[504], lumberyards[504]}), .bottom_left({trees[552], lumberyards[552]}), .bottom({trees[553], lumberyards[553]}), .bottom_right({trees[554], lumberyards[554]}), .init(2'b00), .state({trees[503], lumberyards[503]}));
acre acre_10_4 (.clk(clk), .en(en), .top_left({trees[453], lumberyards[453]}), .top({trees[454], lumberyards[454]}), .top_right({trees[455], lumberyards[455]}), .left({trees[503], lumberyards[503]}), .right({trees[505], lumberyards[505]}), .bottom_left({trees[553], lumberyards[553]}), .bottom({trees[554], lumberyards[554]}), .bottom_right({trees[555], lumberyards[555]}), .init(2'b10), .state({trees[504], lumberyards[504]}));
acre acre_10_5 (.clk(clk), .en(en), .top_left({trees[454], lumberyards[454]}), .top({trees[455], lumberyards[455]}), .top_right({trees[456], lumberyards[456]}), .left({trees[504], lumberyards[504]}), .right({trees[506], lumberyards[506]}), .bottom_left({trees[554], lumberyards[554]}), .bottom({trees[555], lumberyards[555]}), .bottom_right({trees[556], lumberyards[556]}), .init(2'b01), .state({trees[505], lumberyards[505]}));
acre acre_10_6 (.clk(clk), .en(en), .top_left({trees[455], lumberyards[455]}), .top({trees[456], lumberyards[456]}), .top_right({trees[457], lumberyards[457]}), .left({trees[505], lumberyards[505]}), .right({trees[507], lumberyards[507]}), .bottom_left({trees[555], lumberyards[555]}), .bottom({trees[556], lumberyards[556]}), .bottom_right({trees[557], lumberyards[557]}), .init(2'b00), .state({trees[506], lumberyards[506]}));
acre acre_10_7 (.clk(clk), .en(en), .top_left({trees[456], lumberyards[456]}), .top({trees[457], lumberyards[457]}), .top_right({trees[458], lumberyards[458]}), .left({trees[506], lumberyards[506]}), .right({trees[508], lumberyards[508]}), .bottom_left({trees[556], lumberyards[556]}), .bottom({trees[557], lumberyards[557]}), .bottom_right({trees[558], lumberyards[558]}), .init(2'b00), .state({trees[507], lumberyards[507]}));
acre acre_10_8 (.clk(clk), .en(en), .top_left({trees[457], lumberyards[457]}), .top({trees[458], lumberyards[458]}), .top_right({trees[459], lumberyards[459]}), .left({trees[507], lumberyards[507]}), .right({trees[509], lumberyards[509]}), .bottom_left({trees[557], lumberyards[557]}), .bottom({trees[558], lumberyards[558]}), .bottom_right({trees[559], lumberyards[559]}), .init(2'b00), .state({trees[508], lumberyards[508]}));
acre acre_10_9 (.clk(clk), .en(en), .top_left({trees[458], lumberyards[458]}), .top({trees[459], lumberyards[459]}), .top_right({trees[460], lumberyards[460]}), .left({trees[508], lumberyards[508]}), .right({trees[510], lumberyards[510]}), .bottom_left({trees[558], lumberyards[558]}), .bottom({trees[559], lumberyards[559]}), .bottom_right({trees[560], lumberyards[560]}), .init(2'b00), .state({trees[509], lumberyards[509]}));
acre acre_10_10 (.clk(clk), .en(en), .top_left({trees[459], lumberyards[459]}), .top({trees[460], lumberyards[460]}), .top_right({trees[461], lumberyards[461]}), .left({trees[509], lumberyards[509]}), .right({trees[511], lumberyards[511]}), .bottom_left({trees[559], lumberyards[559]}), .bottom({trees[560], lumberyards[560]}), .bottom_right({trees[561], lumberyards[561]}), .init(2'b01), .state({trees[510], lumberyards[510]}));
acre acre_10_11 (.clk(clk), .en(en), .top_left({trees[460], lumberyards[460]}), .top({trees[461], lumberyards[461]}), .top_right({trees[462], lumberyards[462]}), .left({trees[510], lumberyards[510]}), .right({trees[512], lumberyards[512]}), .bottom_left({trees[560], lumberyards[560]}), .bottom({trees[561], lumberyards[561]}), .bottom_right({trees[562], lumberyards[562]}), .init(2'b00), .state({trees[511], lumberyards[511]}));
acre acre_10_12 (.clk(clk), .en(en), .top_left({trees[461], lumberyards[461]}), .top({trees[462], lumberyards[462]}), .top_right({trees[463], lumberyards[463]}), .left({trees[511], lumberyards[511]}), .right({trees[513], lumberyards[513]}), .bottom_left({trees[561], lumberyards[561]}), .bottom({trees[562], lumberyards[562]}), .bottom_right({trees[563], lumberyards[563]}), .init(2'b00), .state({trees[512], lumberyards[512]}));
acre acre_10_13 (.clk(clk), .en(en), .top_left({trees[462], lumberyards[462]}), .top({trees[463], lumberyards[463]}), .top_right({trees[464], lumberyards[464]}), .left({trees[512], lumberyards[512]}), .right({trees[514], lumberyards[514]}), .bottom_left({trees[562], lumberyards[562]}), .bottom({trees[563], lumberyards[563]}), .bottom_right({trees[564], lumberyards[564]}), .init(2'b00), .state({trees[513], lumberyards[513]}));
acre acre_10_14 (.clk(clk), .en(en), .top_left({trees[463], lumberyards[463]}), .top({trees[464], lumberyards[464]}), .top_right({trees[465], lumberyards[465]}), .left({trees[513], lumberyards[513]}), .right({trees[515], lumberyards[515]}), .bottom_left({trees[563], lumberyards[563]}), .bottom({trees[564], lumberyards[564]}), .bottom_right({trees[565], lumberyards[565]}), .init(2'b00), .state({trees[514], lumberyards[514]}));
acre acre_10_15 (.clk(clk), .en(en), .top_left({trees[464], lumberyards[464]}), .top({trees[465], lumberyards[465]}), .top_right({trees[466], lumberyards[466]}), .left({trees[514], lumberyards[514]}), .right({trees[516], lumberyards[516]}), .bottom_left({trees[564], lumberyards[564]}), .bottom({trees[565], lumberyards[565]}), .bottom_right({trees[566], lumberyards[566]}), .init(2'b01), .state({trees[515], lumberyards[515]}));
acre acre_10_16 (.clk(clk), .en(en), .top_left({trees[465], lumberyards[465]}), .top({trees[466], lumberyards[466]}), .top_right({trees[467], lumberyards[467]}), .left({trees[515], lumberyards[515]}), .right({trees[517], lumberyards[517]}), .bottom_left({trees[565], lumberyards[565]}), .bottom({trees[566], lumberyards[566]}), .bottom_right({trees[567], lumberyards[567]}), .init(2'b00), .state({trees[516], lumberyards[516]}));
acre acre_10_17 (.clk(clk), .en(en), .top_left({trees[466], lumberyards[466]}), .top({trees[467], lumberyards[467]}), .top_right({trees[468], lumberyards[468]}), .left({trees[516], lumberyards[516]}), .right({trees[518], lumberyards[518]}), .bottom_left({trees[566], lumberyards[566]}), .bottom({trees[567], lumberyards[567]}), .bottom_right({trees[568], lumberyards[568]}), .init(2'b10), .state({trees[517], lumberyards[517]}));
acre acre_10_18 (.clk(clk), .en(en), .top_left({trees[467], lumberyards[467]}), .top({trees[468], lumberyards[468]}), .top_right({trees[469], lumberyards[469]}), .left({trees[517], lumberyards[517]}), .right({trees[519], lumberyards[519]}), .bottom_left({trees[567], lumberyards[567]}), .bottom({trees[568], lumberyards[568]}), .bottom_right({trees[569], lumberyards[569]}), .init(2'b10), .state({trees[518], lumberyards[518]}));
acre acre_10_19 (.clk(clk), .en(en), .top_left({trees[468], lumberyards[468]}), .top({trees[469], lumberyards[469]}), .top_right({trees[470], lumberyards[470]}), .left({trees[518], lumberyards[518]}), .right({trees[520], lumberyards[520]}), .bottom_left({trees[568], lumberyards[568]}), .bottom({trees[569], lumberyards[569]}), .bottom_right({trees[570], lumberyards[570]}), .init(2'b10), .state({trees[519], lumberyards[519]}));
acre acre_10_20 (.clk(clk), .en(en), .top_left({trees[469], lumberyards[469]}), .top({trees[470], lumberyards[470]}), .top_right({trees[471], lumberyards[471]}), .left({trees[519], lumberyards[519]}), .right({trees[521], lumberyards[521]}), .bottom_left({trees[569], lumberyards[569]}), .bottom({trees[570], lumberyards[570]}), .bottom_right({trees[571], lumberyards[571]}), .init(2'b00), .state({trees[520], lumberyards[520]}));
acre acre_10_21 (.clk(clk), .en(en), .top_left({trees[470], lumberyards[470]}), .top({trees[471], lumberyards[471]}), .top_right({trees[472], lumberyards[472]}), .left({trees[520], lumberyards[520]}), .right({trees[522], lumberyards[522]}), .bottom_left({trees[570], lumberyards[570]}), .bottom({trees[571], lumberyards[571]}), .bottom_right({trees[572], lumberyards[572]}), .init(2'b00), .state({trees[521], lumberyards[521]}));
acre acre_10_22 (.clk(clk), .en(en), .top_left({trees[471], lumberyards[471]}), .top({trees[472], lumberyards[472]}), .top_right({trees[473], lumberyards[473]}), .left({trees[521], lumberyards[521]}), .right({trees[523], lumberyards[523]}), .bottom_left({trees[571], lumberyards[571]}), .bottom({trees[572], lumberyards[572]}), .bottom_right({trees[573], lumberyards[573]}), .init(2'b00), .state({trees[522], lumberyards[522]}));
acre acre_10_23 (.clk(clk), .en(en), .top_left({trees[472], lumberyards[472]}), .top({trees[473], lumberyards[473]}), .top_right({trees[474], lumberyards[474]}), .left({trees[522], lumberyards[522]}), .right({trees[524], lumberyards[524]}), .bottom_left({trees[572], lumberyards[572]}), .bottom({trees[573], lumberyards[573]}), .bottom_right({trees[574], lumberyards[574]}), .init(2'b01), .state({trees[523], lumberyards[523]}));
acre acre_10_24 (.clk(clk), .en(en), .top_left({trees[473], lumberyards[473]}), .top({trees[474], lumberyards[474]}), .top_right({trees[475], lumberyards[475]}), .left({trees[523], lumberyards[523]}), .right({trees[525], lumberyards[525]}), .bottom_left({trees[573], lumberyards[573]}), .bottom({trees[574], lumberyards[574]}), .bottom_right({trees[575], lumberyards[575]}), .init(2'b00), .state({trees[524], lumberyards[524]}));
acre acre_10_25 (.clk(clk), .en(en), .top_left({trees[474], lumberyards[474]}), .top({trees[475], lumberyards[475]}), .top_right({trees[476], lumberyards[476]}), .left({trees[524], lumberyards[524]}), .right({trees[526], lumberyards[526]}), .bottom_left({trees[574], lumberyards[574]}), .bottom({trees[575], lumberyards[575]}), .bottom_right({trees[576], lumberyards[576]}), .init(2'b00), .state({trees[525], lumberyards[525]}));
acre acre_10_26 (.clk(clk), .en(en), .top_left({trees[475], lumberyards[475]}), .top({trees[476], lumberyards[476]}), .top_right({trees[477], lumberyards[477]}), .left({trees[525], lumberyards[525]}), .right({trees[527], lumberyards[527]}), .bottom_left({trees[575], lumberyards[575]}), .bottom({trees[576], lumberyards[576]}), .bottom_right({trees[577], lumberyards[577]}), .init(2'b00), .state({trees[526], lumberyards[526]}));
acre acre_10_27 (.clk(clk), .en(en), .top_left({trees[476], lumberyards[476]}), .top({trees[477], lumberyards[477]}), .top_right({trees[478], lumberyards[478]}), .left({trees[526], lumberyards[526]}), .right({trees[528], lumberyards[528]}), .bottom_left({trees[576], lumberyards[576]}), .bottom({trees[577], lumberyards[577]}), .bottom_right({trees[578], lumberyards[578]}), .init(2'b00), .state({trees[527], lumberyards[527]}));
acre acre_10_28 (.clk(clk), .en(en), .top_left({trees[477], lumberyards[477]}), .top({trees[478], lumberyards[478]}), .top_right({trees[479], lumberyards[479]}), .left({trees[527], lumberyards[527]}), .right({trees[529], lumberyards[529]}), .bottom_left({trees[577], lumberyards[577]}), .bottom({trees[578], lumberyards[578]}), .bottom_right({trees[579], lumberyards[579]}), .init(2'b00), .state({trees[528], lumberyards[528]}));
acre acre_10_29 (.clk(clk), .en(en), .top_left({trees[478], lumberyards[478]}), .top({trees[479], lumberyards[479]}), .top_right({trees[480], lumberyards[480]}), .left({trees[528], lumberyards[528]}), .right({trees[530], lumberyards[530]}), .bottom_left({trees[578], lumberyards[578]}), .bottom({trees[579], lumberyards[579]}), .bottom_right({trees[580], lumberyards[580]}), .init(2'b00), .state({trees[529], lumberyards[529]}));
acre acre_10_30 (.clk(clk), .en(en), .top_left({trees[479], lumberyards[479]}), .top({trees[480], lumberyards[480]}), .top_right({trees[481], lumberyards[481]}), .left({trees[529], lumberyards[529]}), .right({trees[531], lumberyards[531]}), .bottom_left({trees[579], lumberyards[579]}), .bottom({trees[580], lumberyards[580]}), .bottom_right({trees[581], lumberyards[581]}), .init(2'b00), .state({trees[530], lumberyards[530]}));
acre acre_10_31 (.clk(clk), .en(en), .top_left({trees[480], lumberyards[480]}), .top({trees[481], lumberyards[481]}), .top_right({trees[482], lumberyards[482]}), .left({trees[530], lumberyards[530]}), .right({trees[532], lumberyards[532]}), .bottom_left({trees[580], lumberyards[580]}), .bottom({trees[581], lumberyards[581]}), .bottom_right({trees[582], lumberyards[582]}), .init(2'b00), .state({trees[531], lumberyards[531]}));
acre acre_10_32 (.clk(clk), .en(en), .top_left({trees[481], lumberyards[481]}), .top({trees[482], lumberyards[482]}), .top_right({trees[483], lumberyards[483]}), .left({trees[531], lumberyards[531]}), .right({trees[533], lumberyards[533]}), .bottom_left({trees[581], lumberyards[581]}), .bottom({trees[582], lumberyards[582]}), .bottom_right({trees[583], lumberyards[583]}), .init(2'b00), .state({trees[532], lumberyards[532]}));
acre acre_10_33 (.clk(clk), .en(en), .top_left({trees[482], lumberyards[482]}), .top({trees[483], lumberyards[483]}), .top_right({trees[484], lumberyards[484]}), .left({trees[532], lumberyards[532]}), .right({trees[534], lumberyards[534]}), .bottom_left({trees[582], lumberyards[582]}), .bottom({trees[583], lumberyards[583]}), .bottom_right({trees[584], lumberyards[584]}), .init(2'b10), .state({trees[533], lumberyards[533]}));
acre acre_10_34 (.clk(clk), .en(en), .top_left({trees[483], lumberyards[483]}), .top({trees[484], lumberyards[484]}), .top_right({trees[485], lumberyards[485]}), .left({trees[533], lumberyards[533]}), .right({trees[535], lumberyards[535]}), .bottom_left({trees[583], lumberyards[583]}), .bottom({trees[584], lumberyards[584]}), .bottom_right({trees[585], lumberyards[585]}), .init(2'b10), .state({trees[534], lumberyards[534]}));
acre acre_10_35 (.clk(clk), .en(en), .top_left({trees[484], lumberyards[484]}), .top({trees[485], lumberyards[485]}), .top_right({trees[486], lumberyards[486]}), .left({trees[534], lumberyards[534]}), .right({trees[536], lumberyards[536]}), .bottom_left({trees[584], lumberyards[584]}), .bottom({trees[585], lumberyards[585]}), .bottom_right({trees[586], lumberyards[586]}), .init(2'b10), .state({trees[535], lumberyards[535]}));
acre acre_10_36 (.clk(clk), .en(en), .top_left({trees[485], lumberyards[485]}), .top({trees[486], lumberyards[486]}), .top_right({trees[487], lumberyards[487]}), .left({trees[535], lumberyards[535]}), .right({trees[537], lumberyards[537]}), .bottom_left({trees[585], lumberyards[585]}), .bottom({trees[586], lumberyards[586]}), .bottom_right({trees[587], lumberyards[587]}), .init(2'b01), .state({trees[536], lumberyards[536]}));
acre acre_10_37 (.clk(clk), .en(en), .top_left({trees[486], lumberyards[486]}), .top({trees[487], lumberyards[487]}), .top_right({trees[488], lumberyards[488]}), .left({trees[536], lumberyards[536]}), .right({trees[538], lumberyards[538]}), .bottom_left({trees[586], lumberyards[586]}), .bottom({trees[587], lumberyards[587]}), .bottom_right({trees[588], lumberyards[588]}), .init(2'b00), .state({trees[537], lumberyards[537]}));
acre acre_10_38 (.clk(clk), .en(en), .top_left({trees[487], lumberyards[487]}), .top({trees[488], lumberyards[488]}), .top_right({trees[489], lumberyards[489]}), .left({trees[537], lumberyards[537]}), .right({trees[539], lumberyards[539]}), .bottom_left({trees[587], lumberyards[587]}), .bottom({trees[588], lumberyards[588]}), .bottom_right({trees[589], lumberyards[589]}), .init(2'b00), .state({trees[538], lumberyards[538]}));
acre acre_10_39 (.clk(clk), .en(en), .top_left({trees[488], lumberyards[488]}), .top({trees[489], lumberyards[489]}), .top_right({trees[490], lumberyards[490]}), .left({trees[538], lumberyards[538]}), .right({trees[540], lumberyards[540]}), .bottom_left({trees[588], lumberyards[588]}), .bottom({trees[589], lumberyards[589]}), .bottom_right({trees[590], lumberyards[590]}), .init(2'b00), .state({trees[539], lumberyards[539]}));
acre acre_10_40 (.clk(clk), .en(en), .top_left({trees[489], lumberyards[489]}), .top({trees[490], lumberyards[490]}), .top_right({trees[491], lumberyards[491]}), .left({trees[539], lumberyards[539]}), .right({trees[541], lumberyards[541]}), .bottom_left({trees[589], lumberyards[589]}), .bottom({trees[590], lumberyards[590]}), .bottom_right({trees[591], lumberyards[591]}), .init(2'b00), .state({trees[540], lumberyards[540]}));
acre acre_10_41 (.clk(clk), .en(en), .top_left({trees[490], lumberyards[490]}), .top({trees[491], lumberyards[491]}), .top_right({trees[492], lumberyards[492]}), .left({trees[540], lumberyards[540]}), .right({trees[542], lumberyards[542]}), .bottom_left({trees[590], lumberyards[590]}), .bottom({trees[591], lumberyards[591]}), .bottom_right({trees[592], lumberyards[592]}), .init(2'b01), .state({trees[541], lumberyards[541]}));
acre acre_10_42 (.clk(clk), .en(en), .top_left({trees[491], lumberyards[491]}), .top({trees[492], lumberyards[492]}), .top_right({trees[493], lumberyards[493]}), .left({trees[541], lumberyards[541]}), .right({trees[543], lumberyards[543]}), .bottom_left({trees[591], lumberyards[591]}), .bottom({trees[592], lumberyards[592]}), .bottom_right({trees[593], lumberyards[593]}), .init(2'b00), .state({trees[542], lumberyards[542]}));
acre acre_10_43 (.clk(clk), .en(en), .top_left({trees[492], lumberyards[492]}), .top({trees[493], lumberyards[493]}), .top_right({trees[494], lumberyards[494]}), .left({trees[542], lumberyards[542]}), .right({trees[544], lumberyards[544]}), .bottom_left({trees[592], lumberyards[592]}), .bottom({trees[593], lumberyards[593]}), .bottom_right({trees[594], lumberyards[594]}), .init(2'b00), .state({trees[543], lumberyards[543]}));
acre acre_10_44 (.clk(clk), .en(en), .top_left({trees[493], lumberyards[493]}), .top({trees[494], lumberyards[494]}), .top_right({trees[495], lumberyards[495]}), .left({trees[543], lumberyards[543]}), .right({trees[545], lumberyards[545]}), .bottom_left({trees[593], lumberyards[593]}), .bottom({trees[594], lumberyards[594]}), .bottom_right({trees[595], lumberyards[595]}), .init(2'b00), .state({trees[544], lumberyards[544]}));
acre acre_10_45 (.clk(clk), .en(en), .top_left({trees[494], lumberyards[494]}), .top({trees[495], lumberyards[495]}), .top_right({trees[496], lumberyards[496]}), .left({trees[544], lumberyards[544]}), .right({trees[546], lumberyards[546]}), .bottom_left({trees[594], lumberyards[594]}), .bottom({trees[595], lumberyards[595]}), .bottom_right({trees[596], lumberyards[596]}), .init(2'b10), .state({trees[545], lumberyards[545]}));
acre acre_10_46 (.clk(clk), .en(en), .top_left({trees[495], lumberyards[495]}), .top({trees[496], lumberyards[496]}), .top_right({trees[497], lumberyards[497]}), .left({trees[545], lumberyards[545]}), .right({trees[547], lumberyards[547]}), .bottom_left({trees[595], lumberyards[595]}), .bottom({trees[596], lumberyards[596]}), .bottom_right({trees[597], lumberyards[597]}), .init(2'b00), .state({trees[546], lumberyards[546]}));
acre acre_10_47 (.clk(clk), .en(en), .top_left({trees[496], lumberyards[496]}), .top({trees[497], lumberyards[497]}), .top_right({trees[498], lumberyards[498]}), .left({trees[546], lumberyards[546]}), .right({trees[548], lumberyards[548]}), .bottom_left({trees[596], lumberyards[596]}), .bottom({trees[597], lumberyards[597]}), .bottom_right({trees[598], lumberyards[598]}), .init(2'b10), .state({trees[547], lumberyards[547]}));
acre acre_10_48 (.clk(clk), .en(en), .top_left({trees[497], lumberyards[497]}), .top({trees[498], lumberyards[498]}), .top_right({trees[499], lumberyards[499]}), .left({trees[547], lumberyards[547]}), .right({trees[549], lumberyards[549]}), .bottom_left({trees[597], lumberyards[597]}), .bottom({trees[598], lumberyards[598]}), .bottom_right({trees[599], lumberyards[599]}), .init(2'b00), .state({trees[548], lumberyards[548]}));
acre acre_10_49 (.clk(clk), .en(en), .top_left({trees[498], lumberyards[498]}), .top({trees[499], lumberyards[499]}), .top_right(2'b0), .left({trees[548], lumberyards[548]}), .right(2'b0), .bottom_left({trees[598], lumberyards[598]}), .bottom({trees[599], lumberyards[599]}), .bottom_right(2'b0), .init(2'b00), .state({trees[549], lumberyards[549]}));
acre acre_11_0 (.clk(clk), .en(en), .top_left(2'b0), .top({trees[500], lumberyards[500]}), .top_right({trees[501], lumberyards[501]}), .left(2'b0), .right({trees[551], lumberyards[551]}), .bottom_left(2'b0), .bottom({trees[600], lumberyards[600]}), .bottom_right({trees[601], lumberyards[601]}), .init(2'b00), .state({trees[550], lumberyards[550]}));
acre acre_11_1 (.clk(clk), .en(en), .top_left({trees[500], lumberyards[500]}), .top({trees[501], lumberyards[501]}), .top_right({trees[502], lumberyards[502]}), .left({trees[550], lumberyards[550]}), .right({trees[552], lumberyards[552]}), .bottom_left({trees[600], lumberyards[600]}), .bottom({trees[601], lumberyards[601]}), .bottom_right({trees[602], lumberyards[602]}), .init(2'b00), .state({trees[551], lumberyards[551]}));
acre acre_11_2 (.clk(clk), .en(en), .top_left({trees[501], lumberyards[501]}), .top({trees[502], lumberyards[502]}), .top_right({trees[503], lumberyards[503]}), .left({trees[551], lumberyards[551]}), .right({trees[553], lumberyards[553]}), .bottom_left({trees[601], lumberyards[601]}), .bottom({trees[602], lumberyards[602]}), .bottom_right({trees[603], lumberyards[603]}), .init(2'b00), .state({trees[552], lumberyards[552]}));
acre acre_11_3 (.clk(clk), .en(en), .top_left({trees[502], lumberyards[502]}), .top({trees[503], lumberyards[503]}), .top_right({trees[504], lumberyards[504]}), .left({trees[552], lumberyards[552]}), .right({trees[554], lumberyards[554]}), .bottom_left({trees[602], lumberyards[602]}), .bottom({trees[603], lumberyards[603]}), .bottom_right({trees[604], lumberyards[604]}), .init(2'b00), .state({trees[553], lumberyards[553]}));
acre acre_11_4 (.clk(clk), .en(en), .top_left({trees[503], lumberyards[503]}), .top({trees[504], lumberyards[504]}), .top_right({trees[505], lumberyards[505]}), .left({trees[553], lumberyards[553]}), .right({trees[555], lumberyards[555]}), .bottom_left({trees[603], lumberyards[603]}), .bottom({trees[604], lumberyards[604]}), .bottom_right({trees[605], lumberyards[605]}), .init(2'b10), .state({trees[554], lumberyards[554]}));
acre acre_11_5 (.clk(clk), .en(en), .top_left({trees[504], lumberyards[504]}), .top({trees[505], lumberyards[505]}), .top_right({trees[506], lumberyards[506]}), .left({trees[554], lumberyards[554]}), .right({trees[556], lumberyards[556]}), .bottom_left({trees[604], lumberyards[604]}), .bottom({trees[605], lumberyards[605]}), .bottom_right({trees[606], lumberyards[606]}), .init(2'b10), .state({trees[555], lumberyards[555]}));
acre acre_11_6 (.clk(clk), .en(en), .top_left({trees[505], lumberyards[505]}), .top({trees[506], lumberyards[506]}), .top_right({trees[507], lumberyards[507]}), .left({trees[555], lumberyards[555]}), .right({trees[557], lumberyards[557]}), .bottom_left({trees[605], lumberyards[605]}), .bottom({trees[606], lumberyards[606]}), .bottom_right({trees[607], lumberyards[607]}), .init(2'b00), .state({trees[556], lumberyards[556]}));
acre acre_11_7 (.clk(clk), .en(en), .top_left({trees[506], lumberyards[506]}), .top({trees[507], lumberyards[507]}), .top_right({trees[508], lumberyards[508]}), .left({trees[556], lumberyards[556]}), .right({trees[558], lumberyards[558]}), .bottom_left({trees[606], lumberyards[606]}), .bottom({trees[607], lumberyards[607]}), .bottom_right({trees[608], lumberyards[608]}), .init(2'b00), .state({trees[557], lumberyards[557]}));
acre acre_11_8 (.clk(clk), .en(en), .top_left({trees[507], lumberyards[507]}), .top({trees[508], lumberyards[508]}), .top_right({trees[509], lumberyards[509]}), .left({trees[557], lumberyards[557]}), .right({trees[559], lumberyards[559]}), .bottom_left({trees[607], lumberyards[607]}), .bottom({trees[608], lumberyards[608]}), .bottom_right({trees[609], lumberyards[609]}), .init(2'b00), .state({trees[558], lumberyards[558]}));
acre acre_11_9 (.clk(clk), .en(en), .top_left({trees[508], lumberyards[508]}), .top({trees[509], lumberyards[509]}), .top_right({trees[510], lumberyards[510]}), .left({trees[558], lumberyards[558]}), .right({trees[560], lumberyards[560]}), .bottom_left({trees[608], lumberyards[608]}), .bottom({trees[609], lumberyards[609]}), .bottom_right({trees[610], lumberyards[610]}), .init(2'b10), .state({trees[559], lumberyards[559]}));
acre acre_11_10 (.clk(clk), .en(en), .top_left({trees[509], lumberyards[509]}), .top({trees[510], lumberyards[510]}), .top_right({trees[511], lumberyards[511]}), .left({trees[559], lumberyards[559]}), .right({trees[561], lumberyards[561]}), .bottom_left({trees[609], lumberyards[609]}), .bottom({trees[610], lumberyards[610]}), .bottom_right({trees[611], lumberyards[611]}), .init(2'b00), .state({trees[560], lumberyards[560]}));
acre acre_11_11 (.clk(clk), .en(en), .top_left({trees[510], lumberyards[510]}), .top({trees[511], lumberyards[511]}), .top_right({trees[512], lumberyards[512]}), .left({trees[560], lumberyards[560]}), .right({trees[562], lumberyards[562]}), .bottom_left({trees[610], lumberyards[610]}), .bottom({trees[611], lumberyards[611]}), .bottom_right({trees[612], lumberyards[612]}), .init(2'b00), .state({trees[561], lumberyards[561]}));
acre acre_11_12 (.clk(clk), .en(en), .top_left({trees[511], lumberyards[511]}), .top({trees[512], lumberyards[512]}), .top_right({trees[513], lumberyards[513]}), .left({trees[561], lumberyards[561]}), .right({trees[563], lumberyards[563]}), .bottom_left({trees[611], lumberyards[611]}), .bottom({trees[612], lumberyards[612]}), .bottom_right({trees[613], lumberyards[613]}), .init(2'b01), .state({trees[562], lumberyards[562]}));
acre acre_11_13 (.clk(clk), .en(en), .top_left({trees[512], lumberyards[512]}), .top({trees[513], lumberyards[513]}), .top_right({trees[514], lumberyards[514]}), .left({trees[562], lumberyards[562]}), .right({trees[564], lumberyards[564]}), .bottom_left({trees[612], lumberyards[612]}), .bottom({trees[613], lumberyards[613]}), .bottom_right({trees[614], lumberyards[614]}), .init(2'b00), .state({trees[563], lumberyards[563]}));
acre acre_11_14 (.clk(clk), .en(en), .top_left({trees[513], lumberyards[513]}), .top({trees[514], lumberyards[514]}), .top_right({trees[515], lumberyards[515]}), .left({trees[563], lumberyards[563]}), .right({trees[565], lumberyards[565]}), .bottom_left({trees[613], lumberyards[613]}), .bottom({trees[614], lumberyards[614]}), .bottom_right({trees[615], lumberyards[615]}), .init(2'b00), .state({trees[564], lumberyards[564]}));
acre acre_11_15 (.clk(clk), .en(en), .top_left({trees[514], lumberyards[514]}), .top({trees[515], lumberyards[515]}), .top_right({trees[516], lumberyards[516]}), .left({trees[564], lumberyards[564]}), .right({trees[566], lumberyards[566]}), .bottom_left({trees[614], lumberyards[614]}), .bottom({trees[615], lumberyards[615]}), .bottom_right({trees[616], lumberyards[616]}), .init(2'b00), .state({trees[565], lumberyards[565]}));
acre acre_11_16 (.clk(clk), .en(en), .top_left({trees[515], lumberyards[515]}), .top({trees[516], lumberyards[516]}), .top_right({trees[517], lumberyards[517]}), .left({trees[565], lumberyards[565]}), .right({trees[567], lumberyards[567]}), .bottom_left({trees[615], lumberyards[615]}), .bottom({trees[616], lumberyards[616]}), .bottom_right({trees[617], lumberyards[617]}), .init(2'b10), .state({trees[566], lumberyards[566]}));
acre acre_11_17 (.clk(clk), .en(en), .top_left({trees[516], lumberyards[516]}), .top({trees[517], lumberyards[517]}), .top_right({trees[518], lumberyards[518]}), .left({trees[566], lumberyards[566]}), .right({trees[568], lumberyards[568]}), .bottom_left({trees[616], lumberyards[616]}), .bottom({trees[617], lumberyards[617]}), .bottom_right({trees[618], lumberyards[618]}), .init(2'b00), .state({trees[567], lumberyards[567]}));
acre acre_11_18 (.clk(clk), .en(en), .top_left({trees[517], lumberyards[517]}), .top({trees[518], lumberyards[518]}), .top_right({trees[519], lumberyards[519]}), .left({trees[567], lumberyards[567]}), .right({trees[569], lumberyards[569]}), .bottom_left({trees[617], lumberyards[617]}), .bottom({trees[618], lumberyards[618]}), .bottom_right({trees[619], lumberyards[619]}), .init(2'b00), .state({trees[568], lumberyards[568]}));
acre acre_11_19 (.clk(clk), .en(en), .top_left({trees[518], lumberyards[518]}), .top({trees[519], lumberyards[519]}), .top_right({trees[520], lumberyards[520]}), .left({trees[568], lumberyards[568]}), .right({trees[570], lumberyards[570]}), .bottom_left({trees[618], lumberyards[618]}), .bottom({trees[619], lumberyards[619]}), .bottom_right({trees[620], lumberyards[620]}), .init(2'b10), .state({trees[569], lumberyards[569]}));
acre acre_11_20 (.clk(clk), .en(en), .top_left({trees[519], lumberyards[519]}), .top({trees[520], lumberyards[520]}), .top_right({trees[521], lumberyards[521]}), .left({trees[569], lumberyards[569]}), .right({trees[571], lumberyards[571]}), .bottom_left({trees[619], lumberyards[619]}), .bottom({trees[620], lumberyards[620]}), .bottom_right({trees[621], lumberyards[621]}), .init(2'b10), .state({trees[570], lumberyards[570]}));
acre acre_11_21 (.clk(clk), .en(en), .top_left({trees[520], lumberyards[520]}), .top({trees[521], lumberyards[521]}), .top_right({trees[522], lumberyards[522]}), .left({trees[570], lumberyards[570]}), .right({trees[572], lumberyards[572]}), .bottom_left({trees[620], lumberyards[620]}), .bottom({trees[621], lumberyards[621]}), .bottom_right({trees[622], lumberyards[622]}), .init(2'b00), .state({trees[571], lumberyards[571]}));
acre acre_11_22 (.clk(clk), .en(en), .top_left({trees[521], lumberyards[521]}), .top({trees[522], lumberyards[522]}), .top_right({trees[523], lumberyards[523]}), .left({trees[571], lumberyards[571]}), .right({trees[573], lumberyards[573]}), .bottom_left({trees[621], lumberyards[621]}), .bottom({trees[622], lumberyards[622]}), .bottom_right({trees[623], lumberyards[623]}), .init(2'b00), .state({trees[572], lumberyards[572]}));
acre acre_11_23 (.clk(clk), .en(en), .top_left({trees[522], lumberyards[522]}), .top({trees[523], lumberyards[523]}), .top_right({trees[524], lumberyards[524]}), .left({trees[572], lumberyards[572]}), .right({trees[574], lumberyards[574]}), .bottom_left({trees[622], lumberyards[622]}), .bottom({trees[623], lumberyards[623]}), .bottom_right({trees[624], lumberyards[624]}), .init(2'b00), .state({trees[573], lumberyards[573]}));
acre acre_11_24 (.clk(clk), .en(en), .top_left({trees[523], lumberyards[523]}), .top({trees[524], lumberyards[524]}), .top_right({trees[525], lumberyards[525]}), .left({trees[573], lumberyards[573]}), .right({trees[575], lumberyards[575]}), .bottom_left({trees[623], lumberyards[623]}), .bottom({trees[624], lumberyards[624]}), .bottom_right({trees[625], lumberyards[625]}), .init(2'b00), .state({trees[574], lumberyards[574]}));
acre acre_11_25 (.clk(clk), .en(en), .top_left({trees[524], lumberyards[524]}), .top({trees[525], lumberyards[525]}), .top_right({trees[526], lumberyards[526]}), .left({trees[574], lumberyards[574]}), .right({trees[576], lumberyards[576]}), .bottom_left({trees[624], lumberyards[624]}), .bottom({trees[625], lumberyards[625]}), .bottom_right({trees[626], lumberyards[626]}), .init(2'b00), .state({trees[575], lumberyards[575]}));
acre acre_11_26 (.clk(clk), .en(en), .top_left({trees[525], lumberyards[525]}), .top({trees[526], lumberyards[526]}), .top_right({trees[527], lumberyards[527]}), .left({trees[575], lumberyards[575]}), .right({trees[577], lumberyards[577]}), .bottom_left({trees[625], lumberyards[625]}), .bottom({trees[626], lumberyards[626]}), .bottom_right({trees[627], lumberyards[627]}), .init(2'b00), .state({trees[576], lumberyards[576]}));
acre acre_11_27 (.clk(clk), .en(en), .top_left({trees[526], lumberyards[526]}), .top({trees[527], lumberyards[527]}), .top_right({trees[528], lumberyards[528]}), .left({trees[576], lumberyards[576]}), .right({trees[578], lumberyards[578]}), .bottom_left({trees[626], lumberyards[626]}), .bottom({trees[627], lumberyards[627]}), .bottom_right({trees[628], lumberyards[628]}), .init(2'b00), .state({trees[577], lumberyards[577]}));
acre acre_11_28 (.clk(clk), .en(en), .top_left({trees[527], lumberyards[527]}), .top({trees[528], lumberyards[528]}), .top_right({trees[529], lumberyards[529]}), .left({trees[577], lumberyards[577]}), .right({trees[579], lumberyards[579]}), .bottom_left({trees[627], lumberyards[627]}), .bottom({trees[628], lumberyards[628]}), .bottom_right({trees[629], lumberyards[629]}), .init(2'b10), .state({trees[578], lumberyards[578]}));
acre acre_11_29 (.clk(clk), .en(en), .top_left({trees[528], lumberyards[528]}), .top({trees[529], lumberyards[529]}), .top_right({trees[530], lumberyards[530]}), .left({trees[578], lumberyards[578]}), .right({trees[580], lumberyards[580]}), .bottom_left({trees[628], lumberyards[628]}), .bottom({trees[629], lumberyards[629]}), .bottom_right({trees[630], lumberyards[630]}), .init(2'b00), .state({trees[579], lumberyards[579]}));
acre acre_11_30 (.clk(clk), .en(en), .top_left({trees[529], lumberyards[529]}), .top({trees[530], lumberyards[530]}), .top_right({trees[531], lumberyards[531]}), .left({trees[579], lumberyards[579]}), .right({trees[581], lumberyards[581]}), .bottom_left({trees[629], lumberyards[629]}), .bottom({trees[630], lumberyards[630]}), .bottom_right({trees[631], lumberyards[631]}), .init(2'b10), .state({trees[580], lumberyards[580]}));
acre acre_11_31 (.clk(clk), .en(en), .top_left({trees[530], lumberyards[530]}), .top({trees[531], lumberyards[531]}), .top_right({trees[532], lumberyards[532]}), .left({trees[580], lumberyards[580]}), .right({trees[582], lumberyards[582]}), .bottom_left({trees[630], lumberyards[630]}), .bottom({trees[631], lumberyards[631]}), .bottom_right({trees[632], lumberyards[632]}), .init(2'b00), .state({trees[581], lumberyards[581]}));
acre acre_11_32 (.clk(clk), .en(en), .top_left({trees[531], lumberyards[531]}), .top({trees[532], lumberyards[532]}), .top_right({trees[533], lumberyards[533]}), .left({trees[581], lumberyards[581]}), .right({trees[583], lumberyards[583]}), .bottom_left({trees[631], lumberyards[631]}), .bottom({trees[632], lumberyards[632]}), .bottom_right({trees[633], lumberyards[633]}), .init(2'b00), .state({trees[582], lumberyards[582]}));
acre acre_11_33 (.clk(clk), .en(en), .top_left({trees[532], lumberyards[532]}), .top({trees[533], lumberyards[533]}), .top_right({trees[534], lumberyards[534]}), .left({trees[582], lumberyards[582]}), .right({trees[584], lumberyards[584]}), .bottom_left({trees[632], lumberyards[632]}), .bottom({trees[633], lumberyards[633]}), .bottom_right({trees[634], lumberyards[634]}), .init(2'b00), .state({trees[583], lumberyards[583]}));
acre acre_11_34 (.clk(clk), .en(en), .top_left({trees[533], lumberyards[533]}), .top({trees[534], lumberyards[534]}), .top_right({trees[535], lumberyards[535]}), .left({trees[583], lumberyards[583]}), .right({trees[585], lumberyards[585]}), .bottom_left({trees[633], lumberyards[633]}), .bottom({trees[634], lumberyards[634]}), .bottom_right({trees[635], lumberyards[635]}), .init(2'b00), .state({trees[584], lumberyards[584]}));
acre acre_11_35 (.clk(clk), .en(en), .top_left({trees[534], lumberyards[534]}), .top({trees[535], lumberyards[535]}), .top_right({trees[536], lumberyards[536]}), .left({trees[584], lumberyards[584]}), .right({trees[586], lumberyards[586]}), .bottom_left({trees[634], lumberyards[634]}), .bottom({trees[635], lumberyards[635]}), .bottom_right({trees[636], lumberyards[636]}), .init(2'b01), .state({trees[585], lumberyards[585]}));
acre acre_11_36 (.clk(clk), .en(en), .top_left({trees[535], lumberyards[535]}), .top({trees[536], lumberyards[536]}), .top_right({trees[537], lumberyards[537]}), .left({trees[585], lumberyards[585]}), .right({trees[587], lumberyards[587]}), .bottom_left({trees[635], lumberyards[635]}), .bottom({trees[636], lumberyards[636]}), .bottom_right({trees[637], lumberyards[637]}), .init(2'b00), .state({trees[586], lumberyards[586]}));
acre acre_11_37 (.clk(clk), .en(en), .top_left({trees[536], lumberyards[536]}), .top({trees[537], lumberyards[537]}), .top_right({trees[538], lumberyards[538]}), .left({trees[586], lumberyards[586]}), .right({trees[588], lumberyards[588]}), .bottom_left({trees[636], lumberyards[636]}), .bottom({trees[637], lumberyards[637]}), .bottom_right({trees[638], lumberyards[638]}), .init(2'b01), .state({trees[587], lumberyards[587]}));
acre acre_11_38 (.clk(clk), .en(en), .top_left({trees[537], lumberyards[537]}), .top({trees[538], lumberyards[538]}), .top_right({trees[539], lumberyards[539]}), .left({trees[587], lumberyards[587]}), .right({trees[589], lumberyards[589]}), .bottom_left({trees[637], lumberyards[637]}), .bottom({trees[638], lumberyards[638]}), .bottom_right({trees[639], lumberyards[639]}), .init(2'b00), .state({trees[588], lumberyards[588]}));
acre acre_11_39 (.clk(clk), .en(en), .top_left({trees[538], lumberyards[538]}), .top({trees[539], lumberyards[539]}), .top_right({trees[540], lumberyards[540]}), .left({trees[588], lumberyards[588]}), .right({trees[590], lumberyards[590]}), .bottom_left({trees[638], lumberyards[638]}), .bottom({trees[639], lumberyards[639]}), .bottom_right({trees[640], lumberyards[640]}), .init(2'b10), .state({trees[589], lumberyards[589]}));
acre acre_11_40 (.clk(clk), .en(en), .top_left({trees[539], lumberyards[539]}), .top({trees[540], lumberyards[540]}), .top_right({trees[541], lumberyards[541]}), .left({trees[589], lumberyards[589]}), .right({trees[591], lumberyards[591]}), .bottom_left({trees[639], lumberyards[639]}), .bottom({trees[640], lumberyards[640]}), .bottom_right({trees[641], lumberyards[641]}), .init(2'b01), .state({trees[590], lumberyards[590]}));
acre acre_11_41 (.clk(clk), .en(en), .top_left({trees[540], lumberyards[540]}), .top({trees[541], lumberyards[541]}), .top_right({trees[542], lumberyards[542]}), .left({trees[590], lumberyards[590]}), .right({trees[592], lumberyards[592]}), .bottom_left({trees[640], lumberyards[640]}), .bottom({trees[641], lumberyards[641]}), .bottom_right({trees[642], lumberyards[642]}), .init(2'b00), .state({trees[591], lumberyards[591]}));
acre acre_11_42 (.clk(clk), .en(en), .top_left({trees[541], lumberyards[541]}), .top({trees[542], lumberyards[542]}), .top_right({trees[543], lumberyards[543]}), .left({trees[591], lumberyards[591]}), .right({trees[593], lumberyards[593]}), .bottom_left({trees[641], lumberyards[641]}), .bottom({trees[642], lumberyards[642]}), .bottom_right({trees[643], lumberyards[643]}), .init(2'b01), .state({trees[592], lumberyards[592]}));
acre acre_11_43 (.clk(clk), .en(en), .top_left({trees[542], lumberyards[542]}), .top({trees[543], lumberyards[543]}), .top_right({trees[544], lumberyards[544]}), .left({trees[592], lumberyards[592]}), .right({trees[594], lumberyards[594]}), .bottom_left({trees[642], lumberyards[642]}), .bottom({trees[643], lumberyards[643]}), .bottom_right({trees[644], lumberyards[644]}), .init(2'b00), .state({trees[593], lumberyards[593]}));
acre acre_11_44 (.clk(clk), .en(en), .top_left({trees[543], lumberyards[543]}), .top({trees[544], lumberyards[544]}), .top_right({trees[545], lumberyards[545]}), .left({trees[593], lumberyards[593]}), .right({trees[595], lumberyards[595]}), .bottom_left({trees[643], lumberyards[643]}), .bottom({trees[644], lumberyards[644]}), .bottom_right({trees[645], lumberyards[645]}), .init(2'b00), .state({trees[594], lumberyards[594]}));
acre acre_11_45 (.clk(clk), .en(en), .top_left({trees[544], lumberyards[544]}), .top({trees[545], lumberyards[545]}), .top_right({trees[546], lumberyards[546]}), .left({trees[594], lumberyards[594]}), .right({trees[596], lumberyards[596]}), .bottom_left({trees[644], lumberyards[644]}), .bottom({trees[645], lumberyards[645]}), .bottom_right({trees[646], lumberyards[646]}), .init(2'b10), .state({trees[595], lumberyards[595]}));
acre acre_11_46 (.clk(clk), .en(en), .top_left({trees[545], lumberyards[545]}), .top({trees[546], lumberyards[546]}), .top_right({trees[547], lumberyards[547]}), .left({trees[595], lumberyards[595]}), .right({trees[597], lumberyards[597]}), .bottom_left({trees[645], lumberyards[645]}), .bottom({trees[646], lumberyards[646]}), .bottom_right({trees[647], lumberyards[647]}), .init(2'b01), .state({trees[596], lumberyards[596]}));
acre acre_11_47 (.clk(clk), .en(en), .top_left({trees[546], lumberyards[546]}), .top({trees[547], lumberyards[547]}), .top_right({trees[548], lumberyards[548]}), .left({trees[596], lumberyards[596]}), .right({trees[598], lumberyards[598]}), .bottom_left({trees[646], lumberyards[646]}), .bottom({trees[647], lumberyards[647]}), .bottom_right({trees[648], lumberyards[648]}), .init(2'b01), .state({trees[597], lumberyards[597]}));
acre acre_11_48 (.clk(clk), .en(en), .top_left({trees[547], lumberyards[547]}), .top({trees[548], lumberyards[548]}), .top_right({trees[549], lumberyards[549]}), .left({trees[597], lumberyards[597]}), .right({trees[599], lumberyards[599]}), .bottom_left({trees[647], lumberyards[647]}), .bottom({trees[648], lumberyards[648]}), .bottom_right({trees[649], lumberyards[649]}), .init(2'b00), .state({trees[598], lumberyards[598]}));
acre acre_11_49 (.clk(clk), .en(en), .top_left({trees[548], lumberyards[548]}), .top({trees[549], lumberyards[549]}), .top_right(2'b0), .left({trees[598], lumberyards[598]}), .right(2'b0), .bottom_left({trees[648], lumberyards[648]}), .bottom({trees[649], lumberyards[649]}), .bottom_right(2'b0), .init(2'b10), .state({trees[599], lumberyards[599]}));
acre acre_12_0 (.clk(clk), .en(en), .top_left(2'b0), .top({trees[550], lumberyards[550]}), .top_right({trees[551], lumberyards[551]}), .left(2'b0), .right({trees[601], lumberyards[601]}), .bottom_left(2'b0), .bottom({trees[650], lumberyards[650]}), .bottom_right({trees[651], lumberyards[651]}), .init(2'b00), .state({trees[600], lumberyards[600]}));
acre acre_12_1 (.clk(clk), .en(en), .top_left({trees[550], lumberyards[550]}), .top({trees[551], lumberyards[551]}), .top_right({trees[552], lumberyards[552]}), .left({trees[600], lumberyards[600]}), .right({trees[602], lumberyards[602]}), .bottom_left({trees[650], lumberyards[650]}), .bottom({trees[651], lumberyards[651]}), .bottom_right({trees[652], lumberyards[652]}), .init(2'b00), .state({trees[601], lumberyards[601]}));
acre acre_12_2 (.clk(clk), .en(en), .top_left({trees[551], lumberyards[551]}), .top({trees[552], lumberyards[552]}), .top_right({trees[553], lumberyards[553]}), .left({trees[601], lumberyards[601]}), .right({trees[603], lumberyards[603]}), .bottom_left({trees[651], lumberyards[651]}), .bottom({trees[652], lumberyards[652]}), .bottom_right({trees[653], lumberyards[653]}), .init(2'b01), .state({trees[602], lumberyards[602]}));
acre acre_12_3 (.clk(clk), .en(en), .top_left({trees[552], lumberyards[552]}), .top({trees[553], lumberyards[553]}), .top_right({trees[554], lumberyards[554]}), .left({trees[602], lumberyards[602]}), .right({trees[604], lumberyards[604]}), .bottom_left({trees[652], lumberyards[652]}), .bottom({trees[653], lumberyards[653]}), .bottom_right({trees[654], lumberyards[654]}), .init(2'b00), .state({trees[603], lumberyards[603]}));
acre acre_12_4 (.clk(clk), .en(en), .top_left({trees[553], lumberyards[553]}), .top({trees[554], lumberyards[554]}), .top_right({trees[555], lumberyards[555]}), .left({trees[603], lumberyards[603]}), .right({trees[605], lumberyards[605]}), .bottom_left({trees[653], lumberyards[653]}), .bottom({trees[654], lumberyards[654]}), .bottom_right({trees[655], lumberyards[655]}), .init(2'b00), .state({trees[604], lumberyards[604]}));
acre acre_12_5 (.clk(clk), .en(en), .top_left({trees[554], lumberyards[554]}), .top({trees[555], lumberyards[555]}), .top_right({trees[556], lumberyards[556]}), .left({trees[604], lumberyards[604]}), .right({trees[606], lumberyards[606]}), .bottom_left({trees[654], lumberyards[654]}), .bottom({trees[655], lumberyards[655]}), .bottom_right({trees[656], lumberyards[656]}), .init(2'b00), .state({trees[605], lumberyards[605]}));
acre acre_12_6 (.clk(clk), .en(en), .top_left({trees[555], lumberyards[555]}), .top({trees[556], lumberyards[556]}), .top_right({trees[557], lumberyards[557]}), .left({trees[605], lumberyards[605]}), .right({trees[607], lumberyards[607]}), .bottom_left({trees[655], lumberyards[655]}), .bottom({trees[656], lumberyards[656]}), .bottom_right({trees[657], lumberyards[657]}), .init(2'b00), .state({trees[606], lumberyards[606]}));
acre acre_12_7 (.clk(clk), .en(en), .top_left({trees[556], lumberyards[556]}), .top({trees[557], lumberyards[557]}), .top_right({trees[558], lumberyards[558]}), .left({trees[606], lumberyards[606]}), .right({trees[608], lumberyards[608]}), .bottom_left({trees[656], lumberyards[656]}), .bottom({trees[657], lumberyards[657]}), .bottom_right({trees[658], lumberyards[658]}), .init(2'b10), .state({trees[607], lumberyards[607]}));
acre acre_12_8 (.clk(clk), .en(en), .top_left({trees[557], lumberyards[557]}), .top({trees[558], lumberyards[558]}), .top_right({trees[559], lumberyards[559]}), .left({trees[607], lumberyards[607]}), .right({trees[609], lumberyards[609]}), .bottom_left({trees[657], lumberyards[657]}), .bottom({trees[658], lumberyards[658]}), .bottom_right({trees[659], lumberyards[659]}), .init(2'b00), .state({trees[608], lumberyards[608]}));
acre acre_12_9 (.clk(clk), .en(en), .top_left({trees[558], lumberyards[558]}), .top({trees[559], lumberyards[559]}), .top_right({trees[560], lumberyards[560]}), .left({trees[608], lumberyards[608]}), .right({trees[610], lumberyards[610]}), .bottom_left({trees[658], lumberyards[658]}), .bottom({trees[659], lumberyards[659]}), .bottom_right({trees[660], lumberyards[660]}), .init(2'b01), .state({trees[609], lumberyards[609]}));
acre acre_12_10 (.clk(clk), .en(en), .top_left({trees[559], lumberyards[559]}), .top({trees[560], lumberyards[560]}), .top_right({trees[561], lumberyards[561]}), .left({trees[609], lumberyards[609]}), .right({trees[611], lumberyards[611]}), .bottom_left({trees[659], lumberyards[659]}), .bottom({trees[660], lumberyards[660]}), .bottom_right({trees[661], lumberyards[661]}), .init(2'b00), .state({trees[610], lumberyards[610]}));
acre acre_12_11 (.clk(clk), .en(en), .top_left({trees[560], lumberyards[560]}), .top({trees[561], lumberyards[561]}), .top_right({trees[562], lumberyards[562]}), .left({trees[610], lumberyards[610]}), .right({trees[612], lumberyards[612]}), .bottom_left({trees[660], lumberyards[660]}), .bottom({trees[661], lumberyards[661]}), .bottom_right({trees[662], lumberyards[662]}), .init(2'b01), .state({trees[611], lumberyards[611]}));
acre acre_12_12 (.clk(clk), .en(en), .top_left({trees[561], lumberyards[561]}), .top({trees[562], lumberyards[562]}), .top_right({trees[563], lumberyards[563]}), .left({trees[611], lumberyards[611]}), .right({trees[613], lumberyards[613]}), .bottom_left({trees[661], lumberyards[661]}), .bottom({trees[662], lumberyards[662]}), .bottom_right({trees[663], lumberyards[663]}), .init(2'b10), .state({trees[612], lumberyards[612]}));
acre acre_12_13 (.clk(clk), .en(en), .top_left({trees[562], lumberyards[562]}), .top({trees[563], lumberyards[563]}), .top_right({trees[564], lumberyards[564]}), .left({trees[612], lumberyards[612]}), .right({trees[614], lumberyards[614]}), .bottom_left({trees[662], lumberyards[662]}), .bottom({trees[663], lumberyards[663]}), .bottom_right({trees[664], lumberyards[664]}), .init(2'b00), .state({trees[613], lumberyards[613]}));
acre acre_12_14 (.clk(clk), .en(en), .top_left({trees[563], lumberyards[563]}), .top({trees[564], lumberyards[564]}), .top_right({trees[565], lumberyards[565]}), .left({trees[613], lumberyards[613]}), .right({trees[615], lumberyards[615]}), .bottom_left({trees[663], lumberyards[663]}), .bottom({trees[664], lumberyards[664]}), .bottom_right({trees[665], lumberyards[665]}), .init(2'b00), .state({trees[614], lumberyards[614]}));
acre acre_12_15 (.clk(clk), .en(en), .top_left({trees[564], lumberyards[564]}), .top({trees[565], lumberyards[565]}), .top_right({trees[566], lumberyards[566]}), .left({trees[614], lumberyards[614]}), .right({trees[616], lumberyards[616]}), .bottom_left({trees[664], lumberyards[664]}), .bottom({trees[665], lumberyards[665]}), .bottom_right({trees[666], lumberyards[666]}), .init(2'b00), .state({trees[615], lumberyards[615]}));
acre acre_12_16 (.clk(clk), .en(en), .top_left({trees[565], lumberyards[565]}), .top({trees[566], lumberyards[566]}), .top_right({trees[567], lumberyards[567]}), .left({trees[615], lumberyards[615]}), .right({trees[617], lumberyards[617]}), .bottom_left({trees[665], lumberyards[665]}), .bottom({trees[666], lumberyards[666]}), .bottom_right({trees[667], lumberyards[667]}), .init(2'b00), .state({trees[616], lumberyards[616]}));
acre acre_12_17 (.clk(clk), .en(en), .top_left({trees[566], lumberyards[566]}), .top({trees[567], lumberyards[567]}), .top_right({trees[568], lumberyards[568]}), .left({trees[616], lumberyards[616]}), .right({trees[618], lumberyards[618]}), .bottom_left({trees[666], lumberyards[666]}), .bottom({trees[667], lumberyards[667]}), .bottom_right({trees[668], lumberyards[668]}), .init(2'b01), .state({trees[617], lumberyards[617]}));
acre acre_12_18 (.clk(clk), .en(en), .top_left({trees[567], lumberyards[567]}), .top({trees[568], lumberyards[568]}), .top_right({trees[569], lumberyards[569]}), .left({trees[617], lumberyards[617]}), .right({trees[619], lumberyards[619]}), .bottom_left({trees[667], lumberyards[667]}), .bottom({trees[668], lumberyards[668]}), .bottom_right({trees[669], lumberyards[669]}), .init(2'b00), .state({trees[618], lumberyards[618]}));
acre acre_12_19 (.clk(clk), .en(en), .top_left({trees[568], lumberyards[568]}), .top({trees[569], lumberyards[569]}), .top_right({trees[570], lumberyards[570]}), .left({trees[618], lumberyards[618]}), .right({trees[620], lumberyards[620]}), .bottom_left({trees[668], lumberyards[668]}), .bottom({trees[669], lumberyards[669]}), .bottom_right({trees[670], lumberyards[670]}), .init(2'b00), .state({trees[619], lumberyards[619]}));
acre acre_12_20 (.clk(clk), .en(en), .top_left({trees[569], lumberyards[569]}), .top({trees[570], lumberyards[570]}), .top_right({trees[571], lumberyards[571]}), .left({trees[619], lumberyards[619]}), .right({trees[621], lumberyards[621]}), .bottom_left({trees[669], lumberyards[669]}), .bottom({trees[670], lumberyards[670]}), .bottom_right({trees[671], lumberyards[671]}), .init(2'b00), .state({trees[620], lumberyards[620]}));
acre acre_12_21 (.clk(clk), .en(en), .top_left({trees[570], lumberyards[570]}), .top({trees[571], lumberyards[571]}), .top_right({trees[572], lumberyards[572]}), .left({trees[620], lumberyards[620]}), .right({trees[622], lumberyards[622]}), .bottom_left({trees[670], lumberyards[670]}), .bottom({trees[671], lumberyards[671]}), .bottom_right({trees[672], lumberyards[672]}), .init(2'b01), .state({trees[621], lumberyards[621]}));
acre acre_12_22 (.clk(clk), .en(en), .top_left({trees[571], lumberyards[571]}), .top({trees[572], lumberyards[572]}), .top_right({trees[573], lumberyards[573]}), .left({trees[621], lumberyards[621]}), .right({trees[623], lumberyards[623]}), .bottom_left({trees[671], lumberyards[671]}), .bottom({trees[672], lumberyards[672]}), .bottom_right({trees[673], lumberyards[673]}), .init(2'b00), .state({trees[622], lumberyards[622]}));
acre acre_12_23 (.clk(clk), .en(en), .top_left({trees[572], lumberyards[572]}), .top({trees[573], lumberyards[573]}), .top_right({trees[574], lumberyards[574]}), .left({trees[622], lumberyards[622]}), .right({trees[624], lumberyards[624]}), .bottom_left({trees[672], lumberyards[672]}), .bottom({trees[673], lumberyards[673]}), .bottom_right({trees[674], lumberyards[674]}), .init(2'b00), .state({trees[623], lumberyards[623]}));
acre acre_12_24 (.clk(clk), .en(en), .top_left({trees[573], lumberyards[573]}), .top({trees[574], lumberyards[574]}), .top_right({trees[575], lumberyards[575]}), .left({trees[623], lumberyards[623]}), .right({trees[625], lumberyards[625]}), .bottom_left({trees[673], lumberyards[673]}), .bottom({trees[674], lumberyards[674]}), .bottom_right({trees[675], lumberyards[675]}), .init(2'b00), .state({trees[624], lumberyards[624]}));
acre acre_12_25 (.clk(clk), .en(en), .top_left({trees[574], lumberyards[574]}), .top({trees[575], lumberyards[575]}), .top_right({trees[576], lumberyards[576]}), .left({trees[624], lumberyards[624]}), .right({trees[626], lumberyards[626]}), .bottom_left({trees[674], lumberyards[674]}), .bottom({trees[675], lumberyards[675]}), .bottom_right({trees[676], lumberyards[676]}), .init(2'b00), .state({trees[625], lumberyards[625]}));
acre acre_12_26 (.clk(clk), .en(en), .top_left({trees[575], lumberyards[575]}), .top({trees[576], lumberyards[576]}), .top_right({trees[577], lumberyards[577]}), .left({trees[625], lumberyards[625]}), .right({trees[627], lumberyards[627]}), .bottom_left({trees[675], lumberyards[675]}), .bottom({trees[676], lumberyards[676]}), .bottom_right({trees[677], lumberyards[677]}), .init(2'b00), .state({trees[626], lumberyards[626]}));
acre acre_12_27 (.clk(clk), .en(en), .top_left({trees[576], lumberyards[576]}), .top({trees[577], lumberyards[577]}), .top_right({trees[578], lumberyards[578]}), .left({trees[626], lumberyards[626]}), .right({trees[628], lumberyards[628]}), .bottom_left({trees[676], lumberyards[676]}), .bottom({trees[677], lumberyards[677]}), .bottom_right({trees[678], lumberyards[678]}), .init(2'b01), .state({trees[627], lumberyards[627]}));
acre acre_12_28 (.clk(clk), .en(en), .top_left({trees[577], lumberyards[577]}), .top({trees[578], lumberyards[578]}), .top_right({trees[579], lumberyards[579]}), .left({trees[627], lumberyards[627]}), .right({trees[629], lumberyards[629]}), .bottom_left({trees[677], lumberyards[677]}), .bottom({trees[678], lumberyards[678]}), .bottom_right({trees[679], lumberyards[679]}), .init(2'b01), .state({trees[628], lumberyards[628]}));
acre acre_12_29 (.clk(clk), .en(en), .top_left({trees[578], lumberyards[578]}), .top({trees[579], lumberyards[579]}), .top_right({trees[580], lumberyards[580]}), .left({trees[628], lumberyards[628]}), .right({trees[630], lumberyards[630]}), .bottom_left({trees[678], lumberyards[678]}), .bottom({trees[679], lumberyards[679]}), .bottom_right({trees[680], lumberyards[680]}), .init(2'b01), .state({trees[629], lumberyards[629]}));
acre acre_12_30 (.clk(clk), .en(en), .top_left({trees[579], lumberyards[579]}), .top({trees[580], lumberyards[580]}), .top_right({trees[581], lumberyards[581]}), .left({trees[629], lumberyards[629]}), .right({trees[631], lumberyards[631]}), .bottom_left({trees[679], lumberyards[679]}), .bottom({trees[680], lumberyards[680]}), .bottom_right({trees[681], lumberyards[681]}), .init(2'b10), .state({trees[630], lumberyards[630]}));
acre acre_12_31 (.clk(clk), .en(en), .top_left({trees[580], lumberyards[580]}), .top({trees[581], lumberyards[581]}), .top_right({trees[582], lumberyards[582]}), .left({trees[630], lumberyards[630]}), .right({trees[632], lumberyards[632]}), .bottom_left({trees[680], lumberyards[680]}), .bottom({trees[681], lumberyards[681]}), .bottom_right({trees[682], lumberyards[682]}), .init(2'b00), .state({trees[631], lumberyards[631]}));
acre acre_12_32 (.clk(clk), .en(en), .top_left({trees[581], lumberyards[581]}), .top({trees[582], lumberyards[582]}), .top_right({trees[583], lumberyards[583]}), .left({trees[631], lumberyards[631]}), .right({trees[633], lumberyards[633]}), .bottom_left({trees[681], lumberyards[681]}), .bottom({trees[682], lumberyards[682]}), .bottom_right({trees[683], lumberyards[683]}), .init(2'b01), .state({trees[632], lumberyards[632]}));
acre acre_12_33 (.clk(clk), .en(en), .top_left({trees[582], lumberyards[582]}), .top({trees[583], lumberyards[583]}), .top_right({trees[584], lumberyards[584]}), .left({trees[632], lumberyards[632]}), .right({trees[634], lumberyards[634]}), .bottom_left({trees[682], lumberyards[682]}), .bottom({trees[683], lumberyards[683]}), .bottom_right({trees[684], lumberyards[684]}), .init(2'b00), .state({trees[633], lumberyards[633]}));
acre acre_12_34 (.clk(clk), .en(en), .top_left({trees[583], lumberyards[583]}), .top({trees[584], lumberyards[584]}), .top_right({trees[585], lumberyards[585]}), .left({trees[633], lumberyards[633]}), .right({trees[635], lumberyards[635]}), .bottom_left({trees[683], lumberyards[683]}), .bottom({trees[684], lumberyards[684]}), .bottom_right({trees[685], lumberyards[685]}), .init(2'b10), .state({trees[634], lumberyards[634]}));
acre acre_12_35 (.clk(clk), .en(en), .top_left({trees[584], lumberyards[584]}), .top({trees[585], lumberyards[585]}), .top_right({trees[586], lumberyards[586]}), .left({trees[634], lumberyards[634]}), .right({trees[636], lumberyards[636]}), .bottom_left({trees[684], lumberyards[684]}), .bottom({trees[685], lumberyards[685]}), .bottom_right({trees[686], lumberyards[686]}), .init(2'b00), .state({trees[635], lumberyards[635]}));
acre acre_12_36 (.clk(clk), .en(en), .top_left({trees[585], lumberyards[585]}), .top({trees[586], lumberyards[586]}), .top_right({trees[587], lumberyards[587]}), .left({trees[635], lumberyards[635]}), .right({trees[637], lumberyards[637]}), .bottom_left({trees[685], lumberyards[685]}), .bottom({trees[686], lumberyards[686]}), .bottom_right({trees[687], lumberyards[687]}), .init(2'b00), .state({trees[636], lumberyards[636]}));
acre acre_12_37 (.clk(clk), .en(en), .top_left({trees[586], lumberyards[586]}), .top({trees[587], lumberyards[587]}), .top_right({trees[588], lumberyards[588]}), .left({trees[636], lumberyards[636]}), .right({trees[638], lumberyards[638]}), .bottom_left({trees[686], lumberyards[686]}), .bottom({trees[687], lumberyards[687]}), .bottom_right({trees[688], lumberyards[688]}), .init(2'b01), .state({trees[637], lumberyards[637]}));
acre acre_12_38 (.clk(clk), .en(en), .top_left({trees[587], lumberyards[587]}), .top({trees[588], lumberyards[588]}), .top_right({trees[589], lumberyards[589]}), .left({trees[637], lumberyards[637]}), .right({trees[639], lumberyards[639]}), .bottom_left({trees[687], lumberyards[687]}), .bottom({trees[688], lumberyards[688]}), .bottom_right({trees[689], lumberyards[689]}), .init(2'b00), .state({trees[638], lumberyards[638]}));
acre acre_12_39 (.clk(clk), .en(en), .top_left({trees[588], lumberyards[588]}), .top({trees[589], lumberyards[589]}), .top_right({trees[590], lumberyards[590]}), .left({trees[638], lumberyards[638]}), .right({trees[640], lumberyards[640]}), .bottom_left({trees[688], lumberyards[688]}), .bottom({trees[689], lumberyards[689]}), .bottom_right({trees[690], lumberyards[690]}), .init(2'b01), .state({trees[639], lumberyards[639]}));
acre acre_12_40 (.clk(clk), .en(en), .top_left({trees[589], lumberyards[589]}), .top({trees[590], lumberyards[590]}), .top_right({trees[591], lumberyards[591]}), .left({trees[639], lumberyards[639]}), .right({trees[641], lumberyards[641]}), .bottom_left({trees[689], lumberyards[689]}), .bottom({trees[690], lumberyards[690]}), .bottom_right({trees[691], lumberyards[691]}), .init(2'b00), .state({trees[640], lumberyards[640]}));
acre acre_12_41 (.clk(clk), .en(en), .top_left({trees[590], lumberyards[590]}), .top({trees[591], lumberyards[591]}), .top_right({trees[592], lumberyards[592]}), .left({trees[640], lumberyards[640]}), .right({trees[642], lumberyards[642]}), .bottom_left({trees[690], lumberyards[690]}), .bottom({trees[691], lumberyards[691]}), .bottom_right({trees[692], lumberyards[692]}), .init(2'b00), .state({trees[641], lumberyards[641]}));
acre acre_12_42 (.clk(clk), .en(en), .top_left({trees[591], lumberyards[591]}), .top({trees[592], lumberyards[592]}), .top_right({trees[593], lumberyards[593]}), .left({trees[641], lumberyards[641]}), .right({trees[643], lumberyards[643]}), .bottom_left({trees[691], lumberyards[691]}), .bottom({trees[692], lumberyards[692]}), .bottom_right({trees[693], lumberyards[693]}), .init(2'b00), .state({trees[642], lumberyards[642]}));
acre acre_12_43 (.clk(clk), .en(en), .top_left({trees[592], lumberyards[592]}), .top({trees[593], lumberyards[593]}), .top_right({trees[594], lumberyards[594]}), .left({trees[642], lumberyards[642]}), .right({trees[644], lumberyards[644]}), .bottom_left({trees[692], lumberyards[692]}), .bottom({trees[693], lumberyards[693]}), .bottom_right({trees[694], lumberyards[694]}), .init(2'b00), .state({trees[643], lumberyards[643]}));
acre acre_12_44 (.clk(clk), .en(en), .top_left({trees[593], lumberyards[593]}), .top({trees[594], lumberyards[594]}), .top_right({trees[595], lumberyards[595]}), .left({trees[643], lumberyards[643]}), .right({trees[645], lumberyards[645]}), .bottom_left({trees[693], lumberyards[693]}), .bottom({trees[694], lumberyards[694]}), .bottom_right({trees[695], lumberyards[695]}), .init(2'b00), .state({trees[644], lumberyards[644]}));
acre acre_12_45 (.clk(clk), .en(en), .top_left({trees[594], lumberyards[594]}), .top({trees[595], lumberyards[595]}), .top_right({trees[596], lumberyards[596]}), .left({trees[644], lumberyards[644]}), .right({trees[646], lumberyards[646]}), .bottom_left({trees[694], lumberyards[694]}), .bottom({trees[695], lumberyards[695]}), .bottom_right({trees[696], lumberyards[696]}), .init(2'b00), .state({trees[645], lumberyards[645]}));
acre acre_12_46 (.clk(clk), .en(en), .top_left({trees[595], lumberyards[595]}), .top({trees[596], lumberyards[596]}), .top_right({trees[597], lumberyards[597]}), .left({trees[645], lumberyards[645]}), .right({trees[647], lumberyards[647]}), .bottom_left({trees[695], lumberyards[695]}), .bottom({trees[696], lumberyards[696]}), .bottom_right({trees[697], lumberyards[697]}), .init(2'b01), .state({trees[646], lumberyards[646]}));
acre acre_12_47 (.clk(clk), .en(en), .top_left({trees[596], lumberyards[596]}), .top({trees[597], lumberyards[597]}), .top_right({trees[598], lumberyards[598]}), .left({trees[646], lumberyards[646]}), .right({trees[648], lumberyards[648]}), .bottom_left({trees[696], lumberyards[696]}), .bottom({trees[697], lumberyards[697]}), .bottom_right({trees[698], lumberyards[698]}), .init(2'b00), .state({trees[647], lumberyards[647]}));
acre acre_12_48 (.clk(clk), .en(en), .top_left({trees[597], lumberyards[597]}), .top({trees[598], lumberyards[598]}), .top_right({trees[599], lumberyards[599]}), .left({trees[647], lumberyards[647]}), .right({trees[649], lumberyards[649]}), .bottom_left({trees[697], lumberyards[697]}), .bottom({trees[698], lumberyards[698]}), .bottom_right({trees[699], lumberyards[699]}), .init(2'b00), .state({trees[648], lumberyards[648]}));
acre acre_12_49 (.clk(clk), .en(en), .top_left({trees[598], lumberyards[598]}), .top({trees[599], lumberyards[599]}), .top_right(2'b0), .left({trees[648], lumberyards[648]}), .right(2'b0), .bottom_left({trees[698], lumberyards[698]}), .bottom({trees[699], lumberyards[699]}), .bottom_right(2'b0), .init(2'b00), .state({trees[649], lumberyards[649]}));
acre acre_13_0 (.clk(clk), .en(en), .top_left(2'b0), .top({trees[600], lumberyards[600]}), .top_right({trees[601], lumberyards[601]}), .left(2'b0), .right({trees[651], lumberyards[651]}), .bottom_left(2'b0), .bottom({trees[700], lumberyards[700]}), .bottom_right({trees[701], lumberyards[701]}), .init(2'b10), .state({trees[650], lumberyards[650]}));
acre acre_13_1 (.clk(clk), .en(en), .top_left({trees[600], lumberyards[600]}), .top({trees[601], lumberyards[601]}), .top_right({trees[602], lumberyards[602]}), .left({trees[650], lumberyards[650]}), .right({trees[652], lumberyards[652]}), .bottom_left({trees[700], lumberyards[700]}), .bottom({trees[701], lumberyards[701]}), .bottom_right({trees[702], lumberyards[702]}), .init(2'b10), .state({trees[651], lumberyards[651]}));
acre acre_13_2 (.clk(clk), .en(en), .top_left({trees[601], lumberyards[601]}), .top({trees[602], lumberyards[602]}), .top_right({trees[603], lumberyards[603]}), .left({trees[651], lumberyards[651]}), .right({trees[653], lumberyards[653]}), .bottom_left({trees[701], lumberyards[701]}), .bottom({trees[702], lumberyards[702]}), .bottom_right({trees[703], lumberyards[703]}), .init(2'b00), .state({trees[652], lumberyards[652]}));
acre acre_13_3 (.clk(clk), .en(en), .top_left({trees[602], lumberyards[602]}), .top({trees[603], lumberyards[603]}), .top_right({trees[604], lumberyards[604]}), .left({trees[652], lumberyards[652]}), .right({trees[654], lumberyards[654]}), .bottom_left({trees[702], lumberyards[702]}), .bottom({trees[703], lumberyards[703]}), .bottom_right({trees[704], lumberyards[704]}), .init(2'b00), .state({trees[653], lumberyards[653]}));
acre acre_13_4 (.clk(clk), .en(en), .top_left({trees[603], lumberyards[603]}), .top({trees[604], lumberyards[604]}), .top_right({trees[605], lumberyards[605]}), .left({trees[653], lumberyards[653]}), .right({trees[655], lumberyards[655]}), .bottom_left({trees[703], lumberyards[703]}), .bottom({trees[704], lumberyards[704]}), .bottom_right({trees[705], lumberyards[705]}), .init(2'b10), .state({trees[654], lumberyards[654]}));
acre acre_13_5 (.clk(clk), .en(en), .top_left({trees[604], lumberyards[604]}), .top({trees[605], lumberyards[605]}), .top_right({trees[606], lumberyards[606]}), .left({trees[654], lumberyards[654]}), .right({trees[656], lumberyards[656]}), .bottom_left({trees[704], lumberyards[704]}), .bottom({trees[705], lumberyards[705]}), .bottom_right({trees[706], lumberyards[706]}), .init(2'b00), .state({trees[655], lumberyards[655]}));
acre acre_13_6 (.clk(clk), .en(en), .top_left({trees[605], lumberyards[605]}), .top({trees[606], lumberyards[606]}), .top_right({trees[607], lumberyards[607]}), .left({trees[655], lumberyards[655]}), .right({trees[657], lumberyards[657]}), .bottom_left({trees[705], lumberyards[705]}), .bottom({trees[706], lumberyards[706]}), .bottom_right({trees[707], lumberyards[707]}), .init(2'b00), .state({trees[656], lumberyards[656]}));
acre acre_13_7 (.clk(clk), .en(en), .top_left({trees[606], lumberyards[606]}), .top({trees[607], lumberyards[607]}), .top_right({trees[608], lumberyards[608]}), .left({trees[656], lumberyards[656]}), .right({trees[658], lumberyards[658]}), .bottom_left({trees[706], lumberyards[706]}), .bottom({trees[707], lumberyards[707]}), .bottom_right({trees[708], lumberyards[708]}), .init(2'b00), .state({trees[657], lumberyards[657]}));
acre acre_13_8 (.clk(clk), .en(en), .top_left({trees[607], lumberyards[607]}), .top({trees[608], lumberyards[608]}), .top_right({trees[609], lumberyards[609]}), .left({trees[657], lumberyards[657]}), .right({trees[659], lumberyards[659]}), .bottom_left({trees[707], lumberyards[707]}), .bottom({trees[708], lumberyards[708]}), .bottom_right({trees[709], lumberyards[709]}), .init(2'b01), .state({trees[658], lumberyards[658]}));
acre acre_13_9 (.clk(clk), .en(en), .top_left({trees[608], lumberyards[608]}), .top({trees[609], lumberyards[609]}), .top_right({trees[610], lumberyards[610]}), .left({trees[658], lumberyards[658]}), .right({trees[660], lumberyards[660]}), .bottom_left({trees[708], lumberyards[708]}), .bottom({trees[709], lumberyards[709]}), .bottom_right({trees[710], lumberyards[710]}), .init(2'b00), .state({trees[659], lumberyards[659]}));
acre acre_13_10 (.clk(clk), .en(en), .top_left({trees[609], lumberyards[609]}), .top({trees[610], lumberyards[610]}), .top_right({trees[611], lumberyards[611]}), .left({trees[659], lumberyards[659]}), .right({trees[661], lumberyards[661]}), .bottom_left({trees[709], lumberyards[709]}), .bottom({trees[710], lumberyards[710]}), .bottom_right({trees[711], lumberyards[711]}), .init(2'b00), .state({trees[660], lumberyards[660]}));
acre acre_13_11 (.clk(clk), .en(en), .top_left({trees[610], lumberyards[610]}), .top({trees[611], lumberyards[611]}), .top_right({trees[612], lumberyards[612]}), .left({trees[660], lumberyards[660]}), .right({trees[662], lumberyards[662]}), .bottom_left({trees[710], lumberyards[710]}), .bottom({trees[711], lumberyards[711]}), .bottom_right({trees[712], lumberyards[712]}), .init(2'b10), .state({trees[661], lumberyards[661]}));
acre acre_13_12 (.clk(clk), .en(en), .top_left({trees[611], lumberyards[611]}), .top({trees[612], lumberyards[612]}), .top_right({trees[613], lumberyards[613]}), .left({trees[661], lumberyards[661]}), .right({trees[663], lumberyards[663]}), .bottom_left({trees[711], lumberyards[711]}), .bottom({trees[712], lumberyards[712]}), .bottom_right({trees[713], lumberyards[713]}), .init(2'b00), .state({trees[662], lumberyards[662]}));
acre acre_13_13 (.clk(clk), .en(en), .top_left({trees[612], lumberyards[612]}), .top({trees[613], lumberyards[613]}), .top_right({trees[614], lumberyards[614]}), .left({trees[662], lumberyards[662]}), .right({trees[664], lumberyards[664]}), .bottom_left({trees[712], lumberyards[712]}), .bottom({trees[713], lumberyards[713]}), .bottom_right({trees[714], lumberyards[714]}), .init(2'b00), .state({trees[663], lumberyards[663]}));
acre acre_13_14 (.clk(clk), .en(en), .top_left({trees[613], lumberyards[613]}), .top({trees[614], lumberyards[614]}), .top_right({trees[615], lumberyards[615]}), .left({trees[663], lumberyards[663]}), .right({trees[665], lumberyards[665]}), .bottom_left({trees[713], lumberyards[713]}), .bottom({trees[714], lumberyards[714]}), .bottom_right({trees[715], lumberyards[715]}), .init(2'b00), .state({trees[664], lumberyards[664]}));
acre acre_13_15 (.clk(clk), .en(en), .top_left({trees[614], lumberyards[614]}), .top({trees[615], lumberyards[615]}), .top_right({trees[616], lumberyards[616]}), .left({trees[664], lumberyards[664]}), .right({trees[666], lumberyards[666]}), .bottom_left({trees[714], lumberyards[714]}), .bottom({trees[715], lumberyards[715]}), .bottom_right({trees[716], lumberyards[716]}), .init(2'b10), .state({trees[665], lumberyards[665]}));
acre acre_13_16 (.clk(clk), .en(en), .top_left({trees[615], lumberyards[615]}), .top({trees[616], lumberyards[616]}), .top_right({trees[617], lumberyards[617]}), .left({trees[665], lumberyards[665]}), .right({trees[667], lumberyards[667]}), .bottom_left({trees[715], lumberyards[715]}), .bottom({trees[716], lumberyards[716]}), .bottom_right({trees[717], lumberyards[717]}), .init(2'b10), .state({trees[666], lumberyards[666]}));
acre acre_13_17 (.clk(clk), .en(en), .top_left({trees[616], lumberyards[616]}), .top({trees[617], lumberyards[617]}), .top_right({trees[618], lumberyards[618]}), .left({trees[666], lumberyards[666]}), .right({trees[668], lumberyards[668]}), .bottom_left({trees[716], lumberyards[716]}), .bottom({trees[717], lumberyards[717]}), .bottom_right({trees[718], lumberyards[718]}), .init(2'b10), .state({trees[667], lumberyards[667]}));
acre acre_13_18 (.clk(clk), .en(en), .top_left({trees[617], lumberyards[617]}), .top({trees[618], lumberyards[618]}), .top_right({trees[619], lumberyards[619]}), .left({trees[667], lumberyards[667]}), .right({trees[669], lumberyards[669]}), .bottom_left({trees[717], lumberyards[717]}), .bottom({trees[718], lumberyards[718]}), .bottom_right({trees[719], lumberyards[719]}), .init(2'b10), .state({trees[668], lumberyards[668]}));
acre acre_13_19 (.clk(clk), .en(en), .top_left({trees[618], lumberyards[618]}), .top({trees[619], lumberyards[619]}), .top_right({trees[620], lumberyards[620]}), .left({trees[668], lumberyards[668]}), .right({trees[670], lumberyards[670]}), .bottom_left({trees[718], lumberyards[718]}), .bottom({trees[719], lumberyards[719]}), .bottom_right({trees[720], lumberyards[720]}), .init(2'b00), .state({trees[669], lumberyards[669]}));
acre acre_13_20 (.clk(clk), .en(en), .top_left({trees[619], lumberyards[619]}), .top({trees[620], lumberyards[620]}), .top_right({trees[621], lumberyards[621]}), .left({trees[669], lumberyards[669]}), .right({trees[671], lumberyards[671]}), .bottom_left({trees[719], lumberyards[719]}), .bottom({trees[720], lumberyards[720]}), .bottom_right({trees[721], lumberyards[721]}), .init(2'b01), .state({trees[670], lumberyards[670]}));
acre acre_13_21 (.clk(clk), .en(en), .top_left({trees[620], lumberyards[620]}), .top({trees[621], lumberyards[621]}), .top_right({trees[622], lumberyards[622]}), .left({trees[670], lumberyards[670]}), .right({trees[672], lumberyards[672]}), .bottom_left({trees[720], lumberyards[720]}), .bottom({trees[721], lumberyards[721]}), .bottom_right({trees[722], lumberyards[722]}), .init(2'b10), .state({trees[671], lumberyards[671]}));
acre acre_13_22 (.clk(clk), .en(en), .top_left({trees[621], lumberyards[621]}), .top({trees[622], lumberyards[622]}), .top_right({trees[623], lumberyards[623]}), .left({trees[671], lumberyards[671]}), .right({trees[673], lumberyards[673]}), .bottom_left({trees[721], lumberyards[721]}), .bottom({trees[722], lumberyards[722]}), .bottom_right({trees[723], lumberyards[723]}), .init(2'b00), .state({trees[672], lumberyards[672]}));
acre acre_13_23 (.clk(clk), .en(en), .top_left({trees[622], lumberyards[622]}), .top({trees[623], lumberyards[623]}), .top_right({trees[624], lumberyards[624]}), .left({trees[672], lumberyards[672]}), .right({trees[674], lumberyards[674]}), .bottom_left({trees[722], lumberyards[722]}), .bottom({trees[723], lumberyards[723]}), .bottom_right({trees[724], lumberyards[724]}), .init(2'b10), .state({trees[673], lumberyards[673]}));
acre acre_13_24 (.clk(clk), .en(en), .top_left({trees[623], lumberyards[623]}), .top({trees[624], lumberyards[624]}), .top_right({trees[625], lumberyards[625]}), .left({trees[673], lumberyards[673]}), .right({trees[675], lumberyards[675]}), .bottom_left({trees[723], lumberyards[723]}), .bottom({trees[724], lumberyards[724]}), .bottom_right({trees[725], lumberyards[725]}), .init(2'b10), .state({trees[674], lumberyards[674]}));
acre acre_13_25 (.clk(clk), .en(en), .top_left({trees[624], lumberyards[624]}), .top({trees[625], lumberyards[625]}), .top_right({trees[626], lumberyards[626]}), .left({trees[674], lumberyards[674]}), .right({trees[676], lumberyards[676]}), .bottom_left({trees[724], lumberyards[724]}), .bottom({trees[725], lumberyards[725]}), .bottom_right({trees[726], lumberyards[726]}), .init(2'b00), .state({trees[675], lumberyards[675]}));
acre acre_13_26 (.clk(clk), .en(en), .top_left({trees[625], lumberyards[625]}), .top({trees[626], lumberyards[626]}), .top_right({trees[627], lumberyards[627]}), .left({trees[675], lumberyards[675]}), .right({trees[677], lumberyards[677]}), .bottom_left({trees[725], lumberyards[725]}), .bottom({trees[726], lumberyards[726]}), .bottom_right({trees[727], lumberyards[727]}), .init(2'b00), .state({trees[676], lumberyards[676]}));
acre acre_13_27 (.clk(clk), .en(en), .top_left({trees[626], lumberyards[626]}), .top({trees[627], lumberyards[627]}), .top_right({trees[628], lumberyards[628]}), .left({trees[676], lumberyards[676]}), .right({trees[678], lumberyards[678]}), .bottom_left({trees[726], lumberyards[726]}), .bottom({trees[727], lumberyards[727]}), .bottom_right({trees[728], lumberyards[728]}), .init(2'b00), .state({trees[677], lumberyards[677]}));
acre acre_13_28 (.clk(clk), .en(en), .top_left({trees[627], lumberyards[627]}), .top({trees[628], lumberyards[628]}), .top_right({trees[629], lumberyards[629]}), .left({trees[677], lumberyards[677]}), .right({trees[679], lumberyards[679]}), .bottom_left({trees[727], lumberyards[727]}), .bottom({trees[728], lumberyards[728]}), .bottom_right({trees[729], lumberyards[729]}), .init(2'b00), .state({trees[678], lumberyards[678]}));
acre acre_13_29 (.clk(clk), .en(en), .top_left({trees[628], lumberyards[628]}), .top({trees[629], lumberyards[629]}), .top_right({trees[630], lumberyards[630]}), .left({trees[678], lumberyards[678]}), .right({trees[680], lumberyards[680]}), .bottom_left({trees[728], lumberyards[728]}), .bottom({trees[729], lumberyards[729]}), .bottom_right({trees[730], lumberyards[730]}), .init(2'b00), .state({trees[679], lumberyards[679]}));
acre acre_13_30 (.clk(clk), .en(en), .top_left({trees[629], lumberyards[629]}), .top({trees[630], lumberyards[630]}), .top_right({trees[631], lumberyards[631]}), .left({trees[679], lumberyards[679]}), .right({trees[681], lumberyards[681]}), .bottom_left({trees[729], lumberyards[729]}), .bottom({trees[730], lumberyards[730]}), .bottom_right({trees[731], lumberyards[731]}), .init(2'b01), .state({trees[680], lumberyards[680]}));
acre acre_13_31 (.clk(clk), .en(en), .top_left({trees[630], lumberyards[630]}), .top({trees[631], lumberyards[631]}), .top_right({trees[632], lumberyards[632]}), .left({trees[680], lumberyards[680]}), .right({trees[682], lumberyards[682]}), .bottom_left({trees[730], lumberyards[730]}), .bottom({trees[731], lumberyards[731]}), .bottom_right({trees[732], lumberyards[732]}), .init(2'b00), .state({trees[681], lumberyards[681]}));
acre acre_13_32 (.clk(clk), .en(en), .top_left({trees[631], lumberyards[631]}), .top({trees[632], lumberyards[632]}), .top_right({trees[633], lumberyards[633]}), .left({trees[681], lumberyards[681]}), .right({trees[683], lumberyards[683]}), .bottom_left({trees[731], lumberyards[731]}), .bottom({trees[732], lumberyards[732]}), .bottom_right({trees[733], lumberyards[733]}), .init(2'b00), .state({trees[682], lumberyards[682]}));
acre acre_13_33 (.clk(clk), .en(en), .top_left({trees[632], lumberyards[632]}), .top({trees[633], lumberyards[633]}), .top_right({trees[634], lumberyards[634]}), .left({trees[682], lumberyards[682]}), .right({trees[684], lumberyards[684]}), .bottom_left({trees[732], lumberyards[732]}), .bottom({trees[733], lumberyards[733]}), .bottom_right({trees[734], lumberyards[734]}), .init(2'b00), .state({trees[683], lumberyards[683]}));
acre acre_13_34 (.clk(clk), .en(en), .top_left({trees[633], lumberyards[633]}), .top({trees[634], lumberyards[634]}), .top_right({trees[635], lumberyards[635]}), .left({trees[683], lumberyards[683]}), .right({trees[685], lumberyards[685]}), .bottom_left({trees[733], lumberyards[733]}), .bottom({trees[734], lumberyards[734]}), .bottom_right({trees[735], lumberyards[735]}), .init(2'b00), .state({trees[684], lumberyards[684]}));
acre acre_13_35 (.clk(clk), .en(en), .top_left({trees[634], lumberyards[634]}), .top({trees[635], lumberyards[635]}), .top_right({trees[636], lumberyards[636]}), .left({trees[684], lumberyards[684]}), .right({trees[686], lumberyards[686]}), .bottom_left({trees[734], lumberyards[734]}), .bottom({trees[735], lumberyards[735]}), .bottom_right({trees[736], lumberyards[736]}), .init(2'b01), .state({trees[685], lumberyards[685]}));
acre acre_13_36 (.clk(clk), .en(en), .top_left({trees[635], lumberyards[635]}), .top({trees[636], lumberyards[636]}), .top_right({trees[637], lumberyards[637]}), .left({trees[685], lumberyards[685]}), .right({trees[687], lumberyards[687]}), .bottom_left({trees[735], lumberyards[735]}), .bottom({trees[736], lumberyards[736]}), .bottom_right({trees[737], lumberyards[737]}), .init(2'b01), .state({trees[686], lumberyards[686]}));
acre acre_13_37 (.clk(clk), .en(en), .top_left({trees[636], lumberyards[636]}), .top({trees[637], lumberyards[637]}), .top_right({trees[638], lumberyards[638]}), .left({trees[686], lumberyards[686]}), .right({trees[688], lumberyards[688]}), .bottom_left({trees[736], lumberyards[736]}), .bottom({trees[737], lumberyards[737]}), .bottom_right({trees[738], lumberyards[738]}), .init(2'b01), .state({trees[687], lumberyards[687]}));
acre acre_13_38 (.clk(clk), .en(en), .top_left({trees[637], lumberyards[637]}), .top({trees[638], lumberyards[638]}), .top_right({trees[639], lumberyards[639]}), .left({trees[687], lumberyards[687]}), .right({trees[689], lumberyards[689]}), .bottom_left({trees[737], lumberyards[737]}), .bottom({trees[738], lumberyards[738]}), .bottom_right({trees[739], lumberyards[739]}), .init(2'b00), .state({trees[688], lumberyards[688]}));
acre acre_13_39 (.clk(clk), .en(en), .top_left({trees[638], lumberyards[638]}), .top({trees[639], lumberyards[639]}), .top_right({trees[640], lumberyards[640]}), .left({trees[688], lumberyards[688]}), .right({trees[690], lumberyards[690]}), .bottom_left({trees[738], lumberyards[738]}), .bottom({trees[739], lumberyards[739]}), .bottom_right({trees[740], lumberyards[740]}), .init(2'b00), .state({trees[689], lumberyards[689]}));
acre acre_13_40 (.clk(clk), .en(en), .top_left({trees[639], lumberyards[639]}), .top({trees[640], lumberyards[640]}), .top_right({trees[641], lumberyards[641]}), .left({trees[689], lumberyards[689]}), .right({trees[691], lumberyards[691]}), .bottom_left({trees[739], lumberyards[739]}), .bottom({trees[740], lumberyards[740]}), .bottom_right({trees[741], lumberyards[741]}), .init(2'b10), .state({trees[690], lumberyards[690]}));
acre acre_13_41 (.clk(clk), .en(en), .top_left({trees[640], lumberyards[640]}), .top({trees[641], lumberyards[641]}), .top_right({trees[642], lumberyards[642]}), .left({trees[690], lumberyards[690]}), .right({trees[692], lumberyards[692]}), .bottom_left({trees[740], lumberyards[740]}), .bottom({trees[741], lumberyards[741]}), .bottom_right({trees[742], lumberyards[742]}), .init(2'b01), .state({trees[691], lumberyards[691]}));
acre acre_13_42 (.clk(clk), .en(en), .top_left({trees[641], lumberyards[641]}), .top({trees[642], lumberyards[642]}), .top_right({trees[643], lumberyards[643]}), .left({trees[691], lumberyards[691]}), .right({trees[693], lumberyards[693]}), .bottom_left({trees[741], lumberyards[741]}), .bottom({trees[742], lumberyards[742]}), .bottom_right({trees[743], lumberyards[743]}), .init(2'b01), .state({trees[692], lumberyards[692]}));
acre acre_13_43 (.clk(clk), .en(en), .top_left({trees[642], lumberyards[642]}), .top({trees[643], lumberyards[643]}), .top_right({trees[644], lumberyards[644]}), .left({trees[692], lumberyards[692]}), .right({trees[694], lumberyards[694]}), .bottom_left({trees[742], lumberyards[742]}), .bottom({trees[743], lumberyards[743]}), .bottom_right({trees[744], lumberyards[744]}), .init(2'b10), .state({trees[693], lumberyards[693]}));
acre acre_13_44 (.clk(clk), .en(en), .top_left({trees[643], lumberyards[643]}), .top({trees[644], lumberyards[644]}), .top_right({trees[645], lumberyards[645]}), .left({trees[693], lumberyards[693]}), .right({trees[695], lumberyards[695]}), .bottom_left({trees[743], lumberyards[743]}), .bottom({trees[744], lumberyards[744]}), .bottom_right({trees[745], lumberyards[745]}), .init(2'b00), .state({trees[694], lumberyards[694]}));
acre acre_13_45 (.clk(clk), .en(en), .top_left({trees[644], lumberyards[644]}), .top({trees[645], lumberyards[645]}), .top_right({trees[646], lumberyards[646]}), .left({trees[694], lumberyards[694]}), .right({trees[696], lumberyards[696]}), .bottom_left({trees[744], lumberyards[744]}), .bottom({trees[745], lumberyards[745]}), .bottom_right({trees[746], lumberyards[746]}), .init(2'b00), .state({trees[695], lumberyards[695]}));
acre acre_13_46 (.clk(clk), .en(en), .top_left({trees[645], lumberyards[645]}), .top({trees[646], lumberyards[646]}), .top_right({trees[647], lumberyards[647]}), .left({trees[695], lumberyards[695]}), .right({trees[697], lumberyards[697]}), .bottom_left({trees[745], lumberyards[745]}), .bottom({trees[746], lumberyards[746]}), .bottom_right({trees[747], lumberyards[747]}), .init(2'b00), .state({trees[696], lumberyards[696]}));
acre acre_13_47 (.clk(clk), .en(en), .top_left({trees[646], lumberyards[646]}), .top({trees[647], lumberyards[647]}), .top_right({trees[648], lumberyards[648]}), .left({trees[696], lumberyards[696]}), .right({trees[698], lumberyards[698]}), .bottom_left({trees[746], lumberyards[746]}), .bottom({trees[747], lumberyards[747]}), .bottom_right({trees[748], lumberyards[748]}), .init(2'b00), .state({trees[697], lumberyards[697]}));
acre acre_13_48 (.clk(clk), .en(en), .top_left({trees[647], lumberyards[647]}), .top({trees[648], lumberyards[648]}), .top_right({trees[649], lumberyards[649]}), .left({trees[697], lumberyards[697]}), .right({trees[699], lumberyards[699]}), .bottom_left({trees[747], lumberyards[747]}), .bottom({trees[748], lumberyards[748]}), .bottom_right({trees[749], lumberyards[749]}), .init(2'b00), .state({trees[698], lumberyards[698]}));
acre acre_13_49 (.clk(clk), .en(en), .top_left({trees[648], lumberyards[648]}), .top({trees[649], lumberyards[649]}), .top_right(2'b0), .left({trees[698], lumberyards[698]}), .right(2'b0), .bottom_left({trees[748], lumberyards[748]}), .bottom({trees[749], lumberyards[749]}), .bottom_right(2'b0), .init(2'b10), .state({trees[699], lumberyards[699]}));
acre acre_14_0 (.clk(clk), .en(en), .top_left(2'b0), .top({trees[650], lumberyards[650]}), .top_right({trees[651], lumberyards[651]}), .left(2'b0), .right({trees[701], lumberyards[701]}), .bottom_left(2'b0), .bottom({trees[750], lumberyards[750]}), .bottom_right({trees[751], lumberyards[751]}), .init(2'b00), .state({trees[700], lumberyards[700]}));
acre acre_14_1 (.clk(clk), .en(en), .top_left({trees[650], lumberyards[650]}), .top({trees[651], lumberyards[651]}), .top_right({trees[652], lumberyards[652]}), .left({trees[700], lumberyards[700]}), .right({trees[702], lumberyards[702]}), .bottom_left({trees[750], lumberyards[750]}), .bottom({trees[751], lumberyards[751]}), .bottom_right({trees[752], lumberyards[752]}), .init(2'b00), .state({trees[701], lumberyards[701]}));
acre acre_14_2 (.clk(clk), .en(en), .top_left({trees[651], lumberyards[651]}), .top({trees[652], lumberyards[652]}), .top_right({trees[653], lumberyards[653]}), .left({trees[701], lumberyards[701]}), .right({trees[703], lumberyards[703]}), .bottom_left({trees[751], lumberyards[751]}), .bottom({trees[752], lumberyards[752]}), .bottom_right({trees[753], lumberyards[753]}), .init(2'b00), .state({trees[702], lumberyards[702]}));
acre acre_14_3 (.clk(clk), .en(en), .top_left({trees[652], lumberyards[652]}), .top({trees[653], lumberyards[653]}), .top_right({trees[654], lumberyards[654]}), .left({trees[702], lumberyards[702]}), .right({trees[704], lumberyards[704]}), .bottom_left({trees[752], lumberyards[752]}), .bottom({trees[753], lumberyards[753]}), .bottom_right({trees[754], lumberyards[754]}), .init(2'b00), .state({trees[703], lumberyards[703]}));
acre acre_14_4 (.clk(clk), .en(en), .top_left({trees[653], lumberyards[653]}), .top({trees[654], lumberyards[654]}), .top_right({trees[655], lumberyards[655]}), .left({trees[703], lumberyards[703]}), .right({trees[705], lumberyards[705]}), .bottom_left({trees[753], lumberyards[753]}), .bottom({trees[754], lumberyards[754]}), .bottom_right({trees[755], lumberyards[755]}), .init(2'b00), .state({trees[704], lumberyards[704]}));
acre acre_14_5 (.clk(clk), .en(en), .top_left({trees[654], lumberyards[654]}), .top({trees[655], lumberyards[655]}), .top_right({trees[656], lumberyards[656]}), .left({trees[704], lumberyards[704]}), .right({trees[706], lumberyards[706]}), .bottom_left({trees[754], lumberyards[754]}), .bottom({trees[755], lumberyards[755]}), .bottom_right({trees[756], lumberyards[756]}), .init(2'b00), .state({trees[705], lumberyards[705]}));
acre acre_14_6 (.clk(clk), .en(en), .top_left({trees[655], lumberyards[655]}), .top({trees[656], lumberyards[656]}), .top_right({trees[657], lumberyards[657]}), .left({trees[705], lumberyards[705]}), .right({trees[707], lumberyards[707]}), .bottom_left({trees[755], lumberyards[755]}), .bottom({trees[756], lumberyards[756]}), .bottom_right({trees[757], lumberyards[757]}), .init(2'b10), .state({trees[706], lumberyards[706]}));
acre acre_14_7 (.clk(clk), .en(en), .top_left({trees[656], lumberyards[656]}), .top({trees[657], lumberyards[657]}), .top_right({trees[658], lumberyards[658]}), .left({trees[706], lumberyards[706]}), .right({trees[708], lumberyards[708]}), .bottom_left({trees[756], lumberyards[756]}), .bottom({trees[757], lumberyards[757]}), .bottom_right({trees[758], lumberyards[758]}), .init(2'b10), .state({trees[707], lumberyards[707]}));
acre acre_14_8 (.clk(clk), .en(en), .top_left({trees[657], lumberyards[657]}), .top({trees[658], lumberyards[658]}), .top_right({trees[659], lumberyards[659]}), .left({trees[707], lumberyards[707]}), .right({trees[709], lumberyards[709]}), .bottom_left({trees[757], lumberyards[757]}), .bottom({trees[758], lumberyards[758]}), .bottom_right({trees[759], lumberyards[759]}), .init(2'b00), .state({trees[708], lumberyards[708]}));
acre acre_14_9 (.clk(clk), .en(en), .top_left({trees[658], lumberyards[658]}), .top({trees[659], lumberyards[659]}), .top_right({trees[660], lumberyards[660]}), .left({trees[708], lumberyards[708]}), .right({trees[710], lumberyards[710]}), .bottom_left({trees[758], lumberyards[758]}), .bottom({trees[759], lumberyards[759]}), .bottom_right({trees[760], lumberyards[760]}), .init(2'b10), .state({trees[709], lumberyards[709]}));
acre acre_14_10 (.clk(clk), .en(en), .top_left({trees[659], lumberyards[659]}), .top({trees[660], lumberyards[660]}), .top_right({trees[661], lumberyards[661]}), .left({trees[709], lumberyards[709]}), .right({trees[711], lumberyards[711]}), .bottom_left({trees[759], lumberyards[759]}), .bottom({trees[760], lumberyards[760]}), .bottom_right({trees[761], lumberyards[761]}), .init(2'b10), .state({trees[710], lumberyards[710]}));
acre acre_14_11 (.clk(clk), .en(en), .top_left({trees[660], lumberyards[660]}), .top({trees[661], lumberyards[661]}), .top_right({trees[662], lumberyards[662]}), .left({trees[710], lumberyards[710]}), .right({trees[712], lumberyards[712]}), .bottom_left({trees[760], lumberyards[760]}), .bottom({trees[761], lumberyards[761]}), .bottom_right({trees[762], lumberyards[762]}), .init(2'b01), .state({trees[711], lumberyards[711]}));
acre acre_14_12 (.clk(clk), .en(en), .top_left({trees[661], lumberyards[661]}), .top({trees[662], lumberyards[662]}), .top_right({trees[663], lumberyards[663]}), .left({trees[711], lumberyards[711]}), .right({trees[713], lumberyards[713]}), .bottom_left({trees[761], lumberyards[761]}), .bottom({trees[762], lumberyards[762]}), .bottom_right({trees[763], lumberyards[763]}), .init(2'b01), .state({trees[712], lumberyards[712]}));
acre acre_14_13 (.clk(clk), .en(en), .top_left({trees[662], lumberyards[662]}), .top({trees[663], lumberyards[663]}), .top_right({trees[664], lumberyards[664]}), .left({trees[712], lumberyards[712]}), .right({trees[714], lumberyards[714]}), .bottom_left({trees[762], lumberyards[762]}), .bottom({trees[763], lumberyards[763]}), .bottom_right({trees[764], lumberyards[764]}), .init(2'b10), .state({trees[713], lumberyards[713]}));
acre acre_14_14 (.clk(clk), .en(en), .top_left({trees[663], lumberyards[663]}), .top({trees[664], lumberyards[664]}), .top_right({trees[665], lumberyards[665]}), .left({trees[713], lumberyards[713]}), .right({trees[715], lumberyards[715]}), .bottom_left({trees[763], lumberyards[763]}), .bottom({trees[764], lumberyards[764]}), .bottom_right({trees[765], lumberyards[765]}), .init(2'b10), .state({trees[714], lumberyards[714]}));
acre acre_14_15 (.clk(clk), .en(en), .top_left({trees[664], lumberyards[664]}), .top({trees[665], lumberyards[665]}), .top_right({trees[666], lumberyards[666]}), .left({trees[714], lumberyards[714]}), .right({trees[716], lumberyards[716]}), .bottom_left({trees[764], lumberyards[764]}), .bottom({trees[765], lumberyards[765]}), .bottom_right({trees[766], lumberyards[766]}), .init(2'b00), .state({trees[715], lumberyards[715]}));
acre acre_14_16 (.clk(clk), .en(en), .top_left({trees[665], lumberyards[665]}), .top({trees[666], lumberyards[666]}), .top_right({trees[667], lumberyards[667]}), .left({trees[715], lumberyards[715]}), .right({trees[717], lumberyards[717]}), .bottom_left({trees[765], lumberyards[765]}), .bottom({trees[766], lumberyards[766]}), .bottom_right({trees[767], lumberyards[767]}), .init(2'b00), .state({trees[716], lumberyards[716]}));
acre acre_14_17 (.clk(clk), .en(en), .top_left({trees[666], lumberyards[666]}), .top({trees[667], lumberyards[667]}), .top_right({trees[668], lumberyards[668]}), .left({trees[716], lumberyards[716]}), .right({trees[718], lumberyards[718]}), .bottom_left({trees[766], lumberyards[766]}), .bottom({trees[767], lumberyards[767]}), .bottom_right({trees[768], lumberyards[768]}), .init(2'b00), .state({trees[717], lumberyards[717]}));
acre acre_14_18 (.clk(clk), .en(en), .top_left({trees[667], lumberyards[667]}), .top({trees[668], lumberyards[668]}), .top_right({trees[669], lumberyards[669]}), .left({trees[717], lumberyards[717]}), .right({trees[719], lumberyards[719]}), .bottom_left({trees[767], lumberyards[767]}), .bottom({trees[768], lumberyards[768]}), .bottom_right({trees[769], lumberyards[769]}), .init(2'b01), .state({trees[718], lumberyards[718]}));
acre acre_14_19 (.clk(clk), .en(en), .top_left({trees[668], lumberyards[668]}), .top({trees[669], lumberyards[669]}), .top_right({trees[670], lumberyards[670]}), .left({trees[718], lumberyards[718]}), .right({trees[720], lumberyards[720]}), .bottom_left({trees[768], lumberyards[768]}), .bottom({trees[769], lumberyards[769]}), .bottom_right({trees[770], lumberyards[770]}), .init(2'b00), .state({trees[719], lumberyards[719]}));
acre acre_14_20 (.clk(clk), .en(en), .top_left({trees[669], lumberyards[669]}), .top({trees[670], lumberyards[670]}), .top_right({trees[671], lumberyards[671]}), .left({trees[719], lumberyards[719]}), .right({trees[721], lumberyards[721]}), .bottom_left({trees[769], lumberyards[769]}), .bottom({trees[770], lumberyards[770]}), .bottom_right({trees[771], lumberyards[771]}), .init(2'b00), .state({trees[720], lumberyards[720]}));
acre acre_14_21 (.clk(clk), .en(en), .top_left({trees[670], lumberyards[670]}), .top({trees[671], lumberyards[671]}), .top_right({trees[672], lumberyards[672]}), .left({trees[720], lumberyards[720]}), .right({trees[722], lumberyards[722]}), .bottom_left({trees[770], lumberyards[770]}), .bottom({trees[771], lumberyards[771]}), .bottom_right({trees[772], lumberyards[772]}), .init(2'b10), .state({trees[721], lumberyards[721]}));
acre acre_14_22 (.clk(clk), .en(en), .top_left({trees[671], lumberyards[671]}), .top({trees[672], lumberyards[672]}), .top_right({trees[673], lumberyards[673]}), .left({trees[721], lumberyards[721]}), .right({trees[723], lumberyards[723]}), .bottom_left({trees[771], lumberyards[771]}), .bottom({trees[772], lumberyards[772]}), .bottom_right({trees[773], lumberyards[773]}), .init(2'b10), .state({trees[722], lumberyards[722]}));
acre acre_14_23 (.clk(clk), .en(en), .top_left({trees[672], lumberyards[672]}), .top({trees[673], lumberyards[673]}), .top_right({trees[674], lumberyards[674]}), .left({trees[722], lumberyards[722]}), .right({trees[724], lumberyards[724]}), .bottom_left({trees[772], lumberyards[772]}), .bottom({trees[773], lumberyards[773]}), .bottom_right({trees[774], lumberyards[774]}), .init(2'b00), .state({trees[723], lumberyards[723]}));
acre acre_14_24 (.clk(clk), .en(en), .top_left({trees[673], lumberyards[673]}), .top({trees[674], lumberyards[674]}), .top_right({trees[675], lumberyards[675]}), .left({trees[723], lumberyards[723]}), .right({trees[725], lumberyards[725]}), .bottom_left({trees[773], lumberyards[773]}), .bottom({trees[774], lumberyards[774]}), .bottom_right({trees[775], lumberyards[775]}), .init(2'b00), .state({trees[724], lumberyards[724]}));
acre acre_14_25 (.clk(clk), .en(en), .top_left({trees[674], lumberyards[674]}), .top({trees[675], lumberyards[675]}), .top_right({trees[676], lumberyards[676]}), .left({trees[724], lumberyards[724]}), .right({trees[726], lumberyards[726]}), .bottom_left({trees[774], lumberyards[774]}), .bottom({trees[775], lumberyards[775]}), .bottom_right({trees[776], lumberyards[776]}), .init(2'b00), .state({trees[725], lumberyards[725]}));
acre acre_14_26 (.clk(clk), .en(en), .top_left({trees[675], lumberyards[675]}), .top({trees[676], lumberyards[676]}), .top_right({trees[677], lumberyards[677]}), .left({trees[725], lumberyards[725]}), .right({trees[727], lumberyards[727]}), .bottom_left({trees[775], lumberyards[775]}), .bottom({trees[776], lumberyards[776]}), .bottom_right({trees[777], lumberyards[777]}), .init(2'b10), .state({trees[726], lumberyards[726]}));
acre acre_14_27 (.clk(clk), .en(en), .top_left({trees[676], lumberyards[676]}), .top({trees[677], lumberyards[677]}), .top_right({trees[678], lumberyards[678]}), .left({trees[726], lumberyards[726]}), .right({trees[728], lumberyards[728]}), .bottom_left({trees[776], lumberyards[776]}), .bottom({trees[777], lumberyards[777]}), .bottom_right({trees[778], lumberyards[778]}), .init(2'b10), .state({trees[727], lumberyards[727]}));
acre acre_14_28 (.clk(clk), .en(en), .top_left({trees[677], lumberyards[677]}), .top({trees[678], lumberyards[678]}), .top_right({trees[679], lumberyards[679]}), .left({trees[727], lumberyards[727]}), .right({trees[729], lumberyards[729]}), .bottom_left({trees[777], lumberyards[777]}), .bottom({trees[778], lumberyards[778]}), .bottom_right({trees[779], lumberyards[779]}), .init(2'b00), .state({trees[728], lumberyards[728]}));
acre acre_14_29 (.clk(clk), .en(en), .top_left({trees[678], lumberyards[678]}), .top({trees[679], lumberyards[679]}), .top_right({trees[680], lumberyards[680]}), .left({trees[728], lumberyards[728]}), .right({trees[730], lumberyards[730]}), .bottom_left({trees[778], lumberyards[778]}), .bottom({trees[779], lumberyards[779]}), .bottom_right({trees[780], lumberyards[780]}), .init(2'b10), .state({trees[729], lumberyards[729]}));
acre acre_14_30 (.clk(clk), .en(en), .top_left({trees[679], lumberyards[679]}), .top({trees[680], lumberyards[680]}), .top_right({trees[681], lumberyards[681]}), .left({trees[729], lumberyards[729]}), .right({trees[731], lumberyards[731]}), .bottom_left({trees[779], lumberyards[779]}), .bottom({trees[780], lumberyards[780]}), .bottom_right({trees[781], lumberyards[781]}), .init(2'b10), .state({trees[730], lumberyards[730]}));
acre acre_14_31 (.clk(clk), .en(en), .top_left({trees[680], lumberyards[680]}), .top({trees[681], lumberyards[681]}), .top_right({trees[682], lumberyards[682]}), .left({trees[730], lumberyards[730]}), .right({trees[732], lumberyards[732]}), .bottom_left({trees[780], lumberyards[780]}), .bottom({trees[781], lumberyards[781]}), .bottom_right({trees[782], lumberyards[782]}), .init(2'b01), .state({trees[731], lumberyards[731]}));
acre acre_14_32 (.clk(clk), .en(en), .top_left({trees[681], lumberyards[681]}), .top({trees[682], lumberyards[682]}), .top_right({trees[683], lumberyards[683]}), .left({trees[731], lumberyards[731]}), .right({trees[733], lumberyards[733]}), .bottom_left({trees[781], lumberyards[781]}), .bottom({trees[782], lumberyards[782]}), .bottom_right({trees[783], lumberyards[783]}), .init(2'b00), .state({trees[732], lumberyards[732]}));
acre acre_14_33 (.clk(clk), .en(en), .top_left({trees[682], lumberyards[682]}), .top({trees[683], lumberyards[683]}), .top_right({trees[684], lumberyards[684]}), .left({trees[732], lumberyards[732]}), .right({trees[734], lumberyards[734]}), .bottom_left({trees[782], lumberyards[782]}), .bottom({trees[783], lumberyards[783]}), .bottom_right({trees[784], lumberyards[784]}), .init(2'b01), .state({trees[733], lumberyards[733]}));
acre acre_14_34 (.clk(clk), .en(en), .top_left({trees[683], lumberyards[683]}), .top({trees[684], lumberyards[684]}), .top_right({trees[685], lumberyards[685]}), .left({trees[733], lumberyards[733]}), .right({trees[735], lumberyards[735]}), .bottom_left({trees[783], lumberyards[783]}), .bottom({trees[784], lumberyards[784]}), .bottom_right({trees[785], lumberyards[785]}), .init(2'b00), .state({trees[734], lumberyards[734]}));
acre acre_14_35 (.clk(clk), .en(en), .top_left({trees[684], lumberyards[684]}), .top({trees[685], lumberyards[685]}), .top_right({trees[686], lumberyards[686]}), .left({trees[734], lumberyards[734]}), .right({trees[736], lumberyards[736]}), .bottom_left({trees[784], lumberyards[784]}), .bottom({trees[785], lumberyards[785]}), .bottom_right({trees[786], lumberyards[786]}), .init(2'b00), .state({trees[735], lumberyards[735]}));
acre acre_14_36 (.clk(clk), .en(en), .top_left({trees[685], lumberyards[685]}), .top({trees[686], lumberyards[686]}), .top_right({trees[687], lumberyards[687]}), .left({trees[735], lumberyards[735]}), .right({trees[737], lumberyards[737]}), .bottom_left({trees[785], lumberyards[785]}), .bottom({trees[786], lumberyards[786]}), .bottom_right({trees[787], lumberyards[787]}), .init(2'b00), .state({trees[736], lumberyards[736]}));
acre acre_14_37 (.clk(clk), .en(en), .top_left({trees[686], lumberyards[686]}), .top({trees[687], lumberyards[687]}), .top_right({trees[688], lumberyards[688]}), .left({trees[736], lumberyards[736]}), .right({trees[738], lumberyards[738]}), .bottom_left({trees[786], lumberyards[786]}), .bottom({trees[787], lumberyards[787]}), .bottom_right({trees[788], lumberyards[788]}), .init(2'b00), .state({trees[737], lumberyards[737]}));
acre acre_14_38 (.clk(clk), .en(en), .top_left({trees[687], lumberyards[687]}), .top({trees[688], lumberyards[688]}), .top_right({trees[689], lumberyards[689]}), .left({trees[737], lumberyards[737]}), .right({trees[739], lumberyards[739]}), .bottom_left({trees[787], lumberyards[787]}), .bottom({trees[788], lumberyards[788]}), .bottom_right({trees[789], lumberyards[789]}), .init(2'b00), .state({trees[738], lumberyards[738]}));
acre acre_14_39 (.clk(clk), .en(en), .top_left({trees[688], lumberyards[688]}), .top({trees[689], lumberyards[689]}), .top_right({trees[690], lumberyards[690]}), .left({trees[738], lumberyards[738]}), .right({trees[740], lumberyards[740]}), .bottom_left({trees[788], lumberyards[788]}), .bottom({trees[789], lumberyards[789]}), .bottom_right({trees[790], lumberyards[790]}), .init(2'b00), .state({trees[739], lumberyards[739]}));
acre acre_14_40 (.clk(clk), .en(en), .top_left({trees[689], lumberyards[689]}), .top({trees[690], lumberyards[690]}), .top_right({trees[691], lumberyards[691]}), .left({trees[739], lumberyards[739]}), .right({trees[741], lumberyards[741]}), .bottom_left({trees[789], lumberyards[789]}), .bottom({trees[790], lumberyards[790]}), .bottom_right({trees[791], lumberyards[791]}), .init(2'b00), .state({trees[740], lumberyards[740]}));
acre acre_14_41 (.clk(clk), .en(en), .top_left({trees[690], lumberyards[690]}), .top({trees[691], lumberyards[691]}), .top_right({trees[692], lumberyards[692]}), .left({trees[740], lumberyards[740]}), .right({trees[742], lumberyards[742]}), .bottom_left({trees[790], lumberyards[790]}), .bottom({trees[791], lumberyards[791]}), .bottom_right({trees[792], lumberyards[792]}), .init(2'b10), .state({trees[741], lumberyards[741]}));
acre acre_14_42 (.clk(clk), .en(en), .top_left({trees[691], lumberyards[691]}), .top({trees[692], lumberyards[692]}), .top_right({trees[693], lumberyards[693]}), .left({trees[741], lumberyards[741]}), .right({trees[743], lumberyards[743]}), .bottom_left({trees[791], lumberyards[791]}), .bottom({trees[792], lumberyards[792]}), .bottom_right({trees[793], lumberyards[793]}), .init(2'b10), .state({trees[742], lumberyards[742]}));
acre acre_14_43 (.clk(clk), .en(en), .top_left({trees[692], lumberyards[692]}), .top({trees[693], lumberyards[693]}), .top_right({trees[694], lumberyards[694]}), .left({trees[742], lumberyards[742]}), .right({trees[744], lumberyards[744]}), .bottom_left({trees[792], lumberyards[792]}), .bottom({trees[793], lumberyards[793]}), .bottom_right({trees[794], lumberyards[794]}), .init(2'b01), .state({trees[743], lumberyards[743]}));
acre acre_14_44 (.clk(clk), .en(en), .top_left({trees[693], lumberyards[693]}), .top({trees[694], lumberyards[694]}), .top_right({trees[695], lumberyards[695]}), .left({trees[743], lumberyards[743]}), .right({trees[745], lumberyards[745]}), .bottom_left({trees[793], lumberyards[793]}), .bottom({trees[794], lumberyards[794]}), .bottom_right({trees[795], lumberyards[795]}), .init(2'b10), .state({trees[744], lumberyards[744]}));
acre acre_14_45 (.clk(clk), .en(en), .top_left({trees[694], lumberyards[694]}), .top({trees[695], lumberyards[695]}), .top_right({trees[696], lumberyards[696]}), .left({trees[744], lumberyards[744]}), .right({trees[746], lumberyards[746]}), .bottom_left({trees[794], lumberyards[794]}), .bottom({trees[795], lumberyards[795]}), .bottom_right({trees[796], lumberyards[796]}), .init(2'b10), .state({trees[745], lumberyards[745]}));
acre acre_14_46 (.clk(clk), .en(en), .top_left({trees[695], lumberyards[695]}), .top({trees[696], lumberyards[696]}), .top_right({trees[697], lumberyards[697]}), .left({trees[745], lumberyards[745]}), .right({trees[747], lumberyards[747]}), .bottom_left({trees[795], lumberyards[795]}), .bottom({trees[796], lumberyards[796]}), .bottom_right({trees[797], lumberyards[797]}), .init(2'b01), .state({trees[746], lumberyards[746]}));
acre acre_14_47 (.clk(clk), .en(en), .top_left({trees[696], lumberyards[696]}), .top({trees[697], lumberyards[697]}), .top_right({trees[698], lumberyards[698]}), .left({trees[746], lumberyards[746]}), .right({trees[748], lumberyards[748]}), .bottom_left({trees[796], lumberyards[796]}), .bottom({trees[797], lumberyards[797]}), .bottom_right({trees[798], lumberyards[798]}), .init(2'b10), .state({trees[747], lumberyards[747]}));
acre acre_14_48 (.clk(clk), .en(en), .top_left({trees[697], lumberyards[697]}), .top({trees[698], lumberyards[698]}), .top_right({trees[699], lumberyards[699]}), .left({trees[747], lumberyards[747]}), .right({trees[749], lumberyards[749]}), .bottom_left({trees[797], lumberyards[797]}), .bottom({trees[798], lumberyards[798]}), .bottom_right({trees[799], lumberyards[799]}), .init(2'b10), .state({trees[748], lumberyards[748]}));
acre acre_14_49 (.clk(clk), .en(en), .top_left({trees[698], lumberyards[698]}), .top({trees[699], lumberyards[699]}), .top_right(2'b0), .left({trees[748], lumberyards[748]}), .right(2'b0), .bottom_left({trees[798], lumberyards[798]}), .bottom({trees[799], lumberyards[799]}), .bottom_right(2'b0), .init(2'b00), .state({trees[749], lumberyards[749]}));
acre acre_15_0 (.clk(clk), .en(en), .top_left(2'b0), .top({trees[700], lumberyards[700]}), .top_right({trees[701], lumberyards[701]}), .left(2'b0), .right({trees[751], lumberyards[751]}), .bottom_left(2'b0), .bottom({trees[800], lumberyards[800]}), .bottom_right({trees[801], lumberyards[801]}), .init(2'b00), .state({trees[750], lumberyards[750]}));
acre acre_15_1 (.clk(clk), .en(en), .top_left({trees[700], lumberyards[700]}), .top({trees[701], lumberyards[701]}), .top_right({trees[702], lumberyards[702]}), .left({trees[750], lumberyards[750]}), .right({trees[752], lumberyards[752]}), .bottom_left({trees[800], lumberyards[800]}), .bottom({trees[801], lumberyards[801]}), .bottom_right({trees[802], lumberyards[802]}), .init(2'b10), .state({trees[751], lumberyards[751]}));
acre acre_15_2 (.clk(clk), .en(en), .top_left({trees[701], lumberyards[701]}), .top({trees[702], lumberyards[702]}), .top_right({trees[703], lumberyards[703]}), .left({trees[751], lumberyards[751]}), .right({trees[753], lumberyards[753]}), .bottom_left({trees[801], lumberyards[801]}), .bottom({trees[802], lumberyards[802]}), .bottom_right({trees[803], lumberyards[803]}), .init(2'b00), .state({trees[752], lumberyards[752]}));
acre acre_15_3 (.clk(clk), .en(en), .top_left({trees[702], lumberyards[702]}), .top({trees[703], lumberyards[703]}), .top_right({trees[704], lumberyards[704]}), .left({trees[752], lumberyards[752]}), .right({trees[754], lumberyards[754]}), .bottom_left({trees[802], lumberyards[802]}), .bottom({trees[803], lumberyards[803]}), .bottom_right({trees[804], lumberyards[804]}), .init(2'b01), .state({trees[753], lumberyards[753]}));
acre acre_15_4 (.clk(clk), .en(en), .top_left({trees[703], lumberyards[703]}), .top({trees[704], lumberyards[704]}), .top_right({trees[705], lumberyards[705]}), .left({trees[753], lumberyards[753]}), .right({trees[755], lumberyards[755]}), .bottom_left({trees[803], lumberyards[803]}), .bottom({trees[804], lumberyards[804]}), .bottom_right({trees[805], lumberyards[805]}), .init(2'b00), .state({trees[754], lumberyards[754]}));
acre acre_15_5 (.clk(clk), .en(en), .top_left({trees[704], lumberyards[704]}), .top({trees[705], lumberyards[705]}), .top_right({trees[706], lumberyards[706]}), .left({trees[754], lumberyards[754]}), .right({trees[756], lumberyards[756]}), .bottom_left({trees[804], lumberyards[804]}), .bottom({trees[805], lumberyards[805]}), .bottom_right({trees[806], lumberyards[806]}), .init(2'b00), .state({trees[755], lumberyards[755]}));
acre acre_15_6 (.clk(clk), .en(en), .top_left({trees[705], lumberyards[705]}), .top({trees[706], lumberyards[706]}), .top_right({trees[707], lumberyards[707]}), .left({trees[755], lumberyards[755]}), .right({trees[757], lumberyards[757]}), .bottom_left({trees[805], lumberyards[805]}), .bottom({trees[806], lumberyards[806]}), .bottom_right({trees[807], lumberyards[807]}), .init(2'b00), .state({trees[756], lumberyards[756]}));
acre acre_15_7 (.clk(clk), .en(en), .top_left({trees[706], lumberyards[706]}), .top({trees[707], lumberyards[707]}), .top_right({trees[708], lumberyards[708]}), .left({trees[756], lumberyards[756]}), .right({trees[758], lumberyards[758]}), .bottom_left({trees[806], lumberyards[806]}), .bottom({trees[807], lumberyards[807]}), .bottom_right({trees[808], lumberyards[808]}), .init(2'b10), .state({trees[757], lumberyards[757]}));
acre acre_15_8 (.clk(clk), .en(en), .top_left({trees[707], lumberyards[707]}), .top({trees[708], lumberyards[708]}), .top_right({trees[709], lumberyards[709]}), .left({trees[757], lumberyards[757]}), .right({trees[759], lumberyards[759]}), .bottom_left({trees[807], lumberyards[807]}), .bottom({trees[808], lumberyards[808]}), .bottom_right({trees[809], lumberyards[809]}), .init(2'b00), .state({trees[758], lumberyards[758]}));
acre acre_15_9 (.clk(clk), .en(en), .top_left({trees[708], lumberyards[708]}), .top({trees[709], lumberyards[709]}), .top_right({trees[710], lumberyards[710]}), .left({trees[758], lumberyards[758]}), .right({trees[760], lumberyards[760]}), .bottom_left({trees[808], lumberyards[808]}), .bottom({trees[809], lumberyards[809]}), .bottom_right({trees[810], lumberyards[810]}), .init(2'b00), .state({trees[759], lumberyards[759]}));
acre acre_15_10 (.clk(clk), .en(en), .top_left({trees[709], lumberyards[709]}), .top({trees[710], lumberyards[710]}), .top_right({trees[711], lumberyards[711]}), .left({trees[759], lumberyards[759]}), .right({trees[761], lumberyards[761]}), .bottom_left({trees[809], lumberyards[809]}), .bottom({trees[810], lumberyards[810]}), .bottom_right({trees[811], lumberyards[811]}), .init(2'b00), .state({trees[760], lumberyards[760]}));
acre acre_15_11 (.clk(clk), .en(en), .top_left({trees[710], lumberyards[710]}), .top({trees[711], lumberyards[711]}), .top_right({trees[712], lumberyards[712]}), .left({trees[760], lumberyards[760]}), .right({trees[762], lumberyards[762]}), .bottom_left({trees[810], lumberyards[810]}), .bottom({trees[811], lumberyards[811]}), .bottom_right({trees[812], lumberyards[812]}), .init(2'b00), .state({trees[761], lumberyards[761]}));
acre acre_15_12 (.clk(clk), .en(en), .top_left({trees[711], lumberyards[711]}), .top({trees[712], lumberyards[712]}), .top_right({trees[713], lumberyards[713]}), .left({trees[761], lumberyards[761]}), .right({trees[763], lumberyards[763]}), .bottom_left({trees[811], lumberyards[811]}), .bottom({trees[812], lumberyards[812]}), .bottom_right({trees[813], lumberyards[813]}), .init(2'b00), .state({trees[762], lumberyards[762]}));
acre acre_15_13 (.clk(clk), .en(en), .top_left({trees[712], lumberyards[712]}), .top({trees[713], lumberyards[713]}), .top_right({trees[714], lumberyards[714]}), .left({trees[762], lumberyards[762]}), .right({trees[764], lumberyards[764]}), .bottom_left({trees[812], lumberyards[812]}), .bottom({trees[813], lumberyards[813]}), .bottom_right({trees[814], lumberyards[814]}), .init(2'b10), .state({trees[763], lumberyards[763]}));
acre acre_15_14 (.clk(clk), .en(en), .top_left({trees[713], lumberyards[713]}), .top({trees[714], lumberyards[714]}), .top_right({trees[715], lumberyards[715]}), .left({trees[763], lumberyards[763]}), .right({trees[765], lumberyards[765]}), .bottom_left({trees[813], lumberyards[813]}), .bottom({trees[814], lumberyards[814]}), .bottom_right({trees[815], lumberyards[815]}), .init(2'b01), .state({trees[764], lumberyards[764]}));
acre acre_15_15 (.clk(clk), .en(en), .top_left({trees[714], lumberyards[714]}), .top({trees[715], lumberyards[715]}), .top_right({trees[716], lumberyards[716]}), .left({trees[764], lumberyards[764]}), .right({trees[766], lumberyards[766]}), .bottom_left({trees[814], lumberyards[814]}), .bottom({trees[815], lumberyards[815]}), .bottom_right({trees[816], lumberyards[816]}), .init(2'b00), .state({trees[765], lumberyards[765]}));
acre acre_15_16 (.clk(clk), .en(en), .top_left({trees[715], lumberyards[715]}), .top({trees[716], lumberyards[716]}), .top_right({trees[717], lumberyards[717]}), .left({trees[765], lumberyards[765]}), .right({trees[767], lumberyards[767]}), .bottom_left({trees[815], lumberyards[815]}), .bottom({trees[816], lumberyards[816]}), .bottom_right({trees[817], lumberyards[817]}), .init(2'b00), .state({trees[766], lumberyards[766]}));
acre acre_15_17 (.clk(clk), .en(en), .top_left({trees[716], lumberyards[716]}), .top({trees[717], lumberyards[717]}), .top_right({trees[718], lumberyards[718]}), .left({trees[766], lumberyards[766]}), .right({trees[768], lumberyards[768]}), .bottom_left({trees[816], lumberyards[816]}), .bottom({trees[817], lumberyards[817]}), .bottom_right({trees[818], lumberyards[818]}), .init(2'b01), .state({trees[767], lumberyards[767]}));
acre acre_15_18 (.clk(clk), .en(en), .top_left({trees[717], lumberyards[717]}), .top({trees[718], lumberyards[718]}), .top_right({trees[719], lumberyards[719]}), .left({trees[767], lumberyards[767]}), .right({trees[769], lumberyards[769]}), .bottom_left({trees[817], lumberyards[817]}), .bottom({trees[818], lumberyards[818]}), .bottom_right({trees[819], lumberyards[819]}), .init(2'b01), .state({trees[768], lumberyards[768]}));
acre acre_15_19 (.clk(clk), .en(en), .top_left({trees[718], lumberyards[718]}), .top({trees[719], lumberyards[719]}), .top_right({trees[720], lumberyards[720]}), .left({trees[768], lumberyards[768]}), .right({trees[770], lumberyards[770]}), .bottom_left({trees[818], lumberyards[818]}), .bottom({trees[819], lumberyards[819]}), .bottom_right({trees[820], lumberyards[820]}), .init(2'b10), .state({trees[769], lumberyards[769]}));
acre acre_15_20 (.clk(clk), .en(en), .top_left({trees[719], lumberyards[719]}), .top({trees[720], lumberyards[720]}), .top_right({trees[721], lumberyards[721]}), .left({trees[769], lumberyards[769]}), .right({trees[771], lumberyards[771]}), .bottom_left({trees[819], lumberyards[819]}), .bottom({trees[820], lumberyards[820]}), .bottom_right({trees[821], lumberyards[821]}), .init(2'b01), .state({trees[770], lumberyards[770]}));
acre acre_15_21 (.clk(clk), .en(en), .top_left({trees[720], lumberyards[720]}), .top({trees[721], lumberyards[721]}), .top_right({trees[722], lumberyards[722]}), .left({trees[770], lumberyards[770]}), .right({trees[772], lumberyards[772]}), .bottom_left({trees[820], lumberyards[820]}), .bottom({trees[821], lumberyards[821]}), .bottom_right({trees[822], lumberyards[822]}), .init(2'b10), .state({trees[771], lumberyards[771]}));
acre acre_15_22 (.clk(clk), .en(en), .top_left({trees[721], lumberyards[721]}), .top({trees[722], lumberyards[722]}), .top_right({trees[723], lumberyards[723]}), .left({trees[771], lumberyards[771]}), .right({trees[773], lumberyards[773]}), .bottom_left({trees[821], lumberyards[821]}), .bottom({trees[822], lumberyards[822]}), .bottom_right({trees[823], lumberyards[823]}), .init(2'b01), .state({trees[772], lumberyards[772]}));
acre acre_15_23 (.clk(clk), .en(en), .top_left({trees[722], lumberyards[722]}), .top({trees[723], lumberyards[723]}), .top_right({trees[724], lumberyards[724]}), .left({trees[772], lumberyards[772]}), .right({trees[774], lumberyards[774]}), .bottom_left({trees[822], lumberyards[822]}), .bottom({trees[823], lumberyards[823]}), .bottom_right({trees[824], lumberyards[824]}), .init(2'b00), .state({trees[773], lumberyards[773]}));
acre acre_15_24 (.clk(clk), .en(en), .top_left({trees[723], lumberyards[723]}), .top({trees[724], lumberyards[724]}), .top_right({trees[725], lumberyards[725]}), .left({trees[773], lumberyards[773]}), .right({trees[775], lumberyards[775]}), .bottom_left({trees[823], lumberyards[823]}), .bottom({trees[824], lumberyards[824]}), .bottom_right({trees[825], lumberyards[825]}), .init(2'b01), .state({trees[774], lumberyards[774]}));
acre acre_15_25 (.clk(clk), .en(en), .top_left({trees[724], lumberyards[724]}), .top({trees[725], lumberyards[725]}), .top_right({trees[726], lumberyards[726]}), .left({trees[774], lumberyards[774]}), .right({trees[776], lumberyards[776]}), .bottom_left({trees[824], lumberyards[824]}), .bottom({trees[825], lumberyards[825]}), .bottom_right({trees[826], lumberyards[826]}), .init(2'b01), .state({trees[775], lumberyards[775]}));
acre acre_15_26 (.clk(clk), .en(en), .top_left({trees[725], lumberyards[725]}), .top({trees[726], lumberyards[726]}), .top_right({trees[727], lumberyards[727]}), .left({trees[775], lumberyards[775]}), .right({trees[777], lumberyards[777]}), .bottom_left({trees[825], lumberyards[825]}), .bottom({trees[826], lumberyards[826]}), .bottom_right({trees[827], lumberyards[827]}), .init(2'b10), .state({trees[776], lumberyards[776]}));
acre acre_15_27 (.clk(clk), .en(en), .top_left({trees[726], lumberyards[726]}), .top({trees[727], lumberyards[727]}), .top_right({trees[728], lumberyards[728]}), .left({trees[776], lumberyards[776]}), .right({trees[778], lumberyards[778]}), .bottom_left({trees[826], lumberyards[826]}), .bottom({trees[827], lumberyards[827]}), .bottom_right({trees[828], lumberyards[828]}), .init(2'b00), .state({trees[777], lumberyards[777]}));
acre acre_15_28 (.clk(clk), .en(en), .top_left({trees[727], lumberyards[727]}), .top({trees[728], lumberyards[728]}), .top_right({trees[729], lumberyards[729]}), .left({trees[777], lumberyards[777]}), .right({trees[779], lumberyards[779]}), .bottom_left({trees[827], lumberyards[827]}), .bottom({trees[828], lumberyards[828]}), .bottom_right({trees[829], lumberyards[829]}), .init(2'b00), .state({trees[778], lumberyards[778]}));
acre acre_15_29 (.clk(clk), .en(en), .top_left({trees[728], lumberyards[728]}), .top({trees[729], lumberyards[729]}), .top_right({trees[730], lumberyards[730]}), .left({trees[778], lumberyards[778]}), .right({trees[780], lumberyards[780]}), .bottom_left({trees[828], lumberyards[828]}), .bottom({trees[829], lumberyards[829]}), .bottom_right({trees[830], lumberyards[830]}), .init(2'b10), .state({trees[779], lumberyards[779]}));
acre acre_15_30 (.clk(clk), .en(en), .top_left({trees[729], lumberyards[729]}), .top({trees[730], lumberyards[730]}), .top_right({trees[731], lumberyards[731]}), .left({trees[779], lumberyards[779]}), .right({trees[781], lumberyards[781]}), .bottom_left({trees[829], lumberyards[829]}), .bottom({trees[830], lumberyards[830]}), .bottom_right({trees[831], lumberyards[831]}), .init(2'b01), .state({trees[780], lumberyards[780]}));
acre acre_15_31 (.clk(clk), .en(en), .top_left({trees[730], lumberyards[730]}), .top({trees[731], lumberyards[731]}), .top_right({trees[732], lumberyards[732]}), .left({trees[780], lumberyards[780]}), .right({trees[782], lumberyards[782]}), .bottom_left({trees[830], lumberyards[830]}), .bottom({trees[831], lumberyards[831]}), .bottom_right({trees[832], lumberyards[832]}), .init(2'b01), .state({trees[781], lumberyards[781]}));
acre acre_15_32 (.clk(clk), .en(en), .top_left({trees[731], lumberyards[731]}), .top({trees[732], lumberyards[732]}), .top_right({trees[733], lumberyards[733]}), .left({trees[781], lumberyards[781]}), .right({trees[783], lumberyards[783]}), .bottom_left({trees[831], lumberyards[831]}), .bottom({trees[832], lumberyards[832]}), .bottom_right({trees[833], lumberyards[833]}), .init(2'b00), .state({trees[782], lumberyards[782]}));
acre acre_15_33 (.clk(clk), .en(en), .top_left({trees[732], lumberyards[732]}), .top({trees[733], lumberyards[733]}), .top_right({trees[734], lumberyards[734]}), .left({trees[782], lumberyards[782]}), .right({trees[784], lumberyards[784]}), .bottom_left({trees[832], lumberyards[832]}), .bottom({trees[833], lumberyards[833]}), .bottom_right({trees[834], lumberyards[834]}), .init(2'b00), .state({trees[783], lumberyards[783]}));
acre acre_15_34 (.clk(clk), .en(en), .top_left({trees[733], lumberyards[733]}), .top({trees[734], lumberyards[734]}), .top_right({trees[735], lumberyards[735]}), .left({trees[783], lumberyards[783]}), .right({trees[785], lumberyards[785]}), .bottom_left({trees[833], lumberyards[833]}), .bottom({trees[834], lumberyards[834]}), .bottom_right({trees[835], lumberyards[835]}), .init(2'b00), .state({trees[784], lumberyards[784]}));
acre acre_15_35 (.clk(clk), .en(en), .top_left({trees[734], lumberyards[734]}), .top({trees[735], lumberyards[735]}), .top_right({trees[736], lumberyards[736]}), .left({trees[784], lumberyards[784]}), .right({trees[786], lumberyards[786]}), .bottom_left({trees[834], lumberyards[834]}), .bottom({trees[835], lumberyards[835]}), .bottom_right({trees[836], lumberyards[836]}), .init(2'b01), .state({trees[785], lumberyards[785]}));
acre acre_15_36 (.clk(clk), .en(en), .top_left({trees[735], lumberyards[735]}), .top({trees[736], lumberyards[736]}), .top_right({trees[737], lumberyards[737]}), .left({trees[785], lumberyards[785]}), .right({trees[787], lumberyards[787]}), .bottom_left({trees[835], lumberyards[835]}), .bottom({trees[836], lumberyards[836]}), .bottom_right({trees[837], lumberyards[837]}), .init(2'b00), .state({trees[786], lumberyards[786]}));
acre acre_15_37 (.clk(clk), .en(en), .top_left({trees[736], lumberyards[736]}), .top({trees[737], lumberyards[737]}), .top_right({trees[738], lumberyards[738]}), .left({trees[786], lumberyards[786]}), .right({trees[788], lumberyards[788]}), .bottom_left({trees[836], lumberyards[836]}), .bottom({trees[837], lumberyards[837]}), .bottom_right({trees[838], lumberyards[838]}), .init(2'b00), .state({trees[787], lumberyards[787]}));
acre acre_15_38 (.clk(clk), .en(en), .top_left({trees[737], lumberyards[737]}), .top({trees[738], lumberyards[738]}), .top_right({trees[739], lumberyards[739]}), .left({trees[787], lumberyards[787]}), .right({trees[789], lumberyards[789]}), .bottom_left({trees[837], lumberyards[837]}), .bottom({trees[838], lumberyards[838]}), .bottom_right({trees[839], lumberyards[839]}), .init(2'b00), .state({trees[788], lumberyards[788]}));
acre acre_15_39 (.clk(clk), .en(en), .top_left({trees[738], lumberyards[738]}), .top({trees[739], lumberyards[739]}), .top_right({trees[740], lumberyards[740]}), .left({trees[788], lumberyards[788]}), .right({trees[790], lumberyards[790]}), .bottom_left({trees[838], lumberyards[838]}), .bottom({trees[839], lumberyards[839]}), .bottom_right({trees[840], lumberyards[840]}), .init(2'b10), .state({trees[789], lumberyards[789]}));
acre acre_15_40 (.clk(clk), .en(en), .top_left({trees[739], lumberyards[739]}), .top({trees[740], lumberyards[740]}), .top_right({trees[741], lumberyards[741]}), .left({trees[789], lumberyards[789]}), .right({trees[791], lumberyards[791]}), .bottom_left({trees[839], lumberyards[839]}), .bottom({trees[840], lumberyards[840]}), .bottom_right({trees[841], lumberyards[841]}), .init(2'b00), .state({trees[790], lumberyards[790]}));
acre acre_15_41 (.clk(clk), .en(en), .top_left({trees[740], lumberyards[740]}), .top({trees[741], lumberyards[741]}), .top_right({trees[742], lumberyards[742]}), .left({trees[790], lumberyards[790]}), .right({trees[792], lumberyards[792]}), .bottom_left({trees[840], lumberyards[840]}), .bottom({trees[841], lumberyards[841]}), .bottom_right({trees[842], lumberyards[842]}), .init(2'b00), .state({trees[791], lumberyards[791]}));
acre acre_15_42 (.clk(clk), .en(en), .top_left({trees[741], lumberyards[741]}), .top({trees[742], lumberyards[742]}), .top_right({trees[743], lumberyards[743]}), .left({trees[791], lumberyards[791]}), .right({trees[793], lumberyards[793]}), .bottom_left({trees[841], lumberyards[841]}), .bottom({trees[842], lumberyards[842]}), .bottom_right({trees[843], lumberyards[843]}), .init(2'b01), .state({trees[792], lumberyards[792]}));
acre acre_15_43 (.clk(clk), .en(en), .top_left({trees[742], lumberyards[742]}), .top({trees[743], lumberyards[743]}), .top_right({trees[744], lumberyards[744]}), .left({trees[792], lumberyards[792]}), .right({trees[794], lumberyards[794]}), .bottom_left({trees[842], lumberyards[842]}), .bottom({trees[843], lumberyards[843]}), .bottom_right({trees[844], lumberyards[844]}), .init(2'b10), .state({trees[793], lumberyards[793]}));
acre acre_15_44 (.clk(clk), .en(en), .top_left({trees[743], lumberyards[743]}), .top({trees[744], lumberyards[744]}), .top_right({trees[745], lumberyards[745]}), .left({trees[793], lumberyards[793]}), .right({trees[795], lumberyards[795]}), .bottom_left({trees[843], lumberyards[843]}), .bottom({trees[844], lumberyards[844]}), .bottom_right({trees[845], lumberyards[845]}), .init(2'b01), .state({trees[794], lumberyards[794]}));
acre acre_15_45 (.clk(clk), .en(en), .top_left({trees[744], lumberyards[744]}), .top({trees[745], lumberyards[745]}), .top_right({trees[746], lumberyards[746]}), .left({trees[794], lumberyards[794]}), .right({trees[796], lumberyards[796]}), .bottom_left({trees[844], lumberyards[844]}), .bottom({trees[845], lumberyards[845]}), .bottom_right({trees[846], lumberyards[846]}), .init(2'b01), .state({trees[795], lumberyards[795]}));
acre acre_15_46 (.clk(clk), .en(en), .top_left({trees[745], lumberyards[745]}), .top({trees[746], lumberyards[746]}), .top_right({trees[747], lumberyards[747]}), .left({trees[795], lumberyards[795]}), .right({trees[797], lumberyards[797]}), .bottom_left({trees[845], lumberyards[845]}), .bottom({trees[846], lumberyards[846]}), .bottom_right({trees[847], lumberyards[847]}), .init(2'b00), .state({trees[796], lumberyards[796]}));
acre acre_15_47 (.clk(clk), .en(en), .top_left({trees[746], lumberyards[746]}), .top({trees[747], lumberyards[747]}), .top_right({trees[748], lumberyards[748]}), .left({trees[796], lumberyards[796]}), .right({trees[798], lumberyards[798]}), .bottom_left({trees[846], lumberyards[846]}), .bottom({trees[847], lumberyards[847]}), .bottom_right({trees[848], lumberyards[848]}), .init(2'b00), .state({trees[797], lumberyards[797]}));
acre acre_15_48 (.clk(clk), .en(en), .top_left({trees[747], lumberyards[747]}), .top({trees[748], lumberyards[748]}), .top_right({trees[749], lumberyards[749]}), .left({trees[797], lumberyards[797]}), .right({trees[799], lumberyards[799]}), .bottom_left({trees[847], lumberyards[847]}), .bottom({trees[848], lumberyards[848]}), .bottom_right({trees[849], lumberyards[849]}), .init(2'b10), .state({trees[798], lumberyards[798]}));
acre acre_15_49 (.clk(clk), .en(en), .top_left({trees[748], lumberyards[748]}), .top({trees[749], lumberyards[749]}), .top_right(2'b0), .left({trees[798], lumberyards[798]}), .right(2'b0), .bottom_left({trees[848], lumberyards[848]}), .bottom({trees[849], lumberyards[849]}), .bottom_right(2'b0), .init(2'b00), .state({trees[799], lumberyards[799]}));
acre acre_16_0 (.clk(clk), .en(en), .top_left(2'b0), .top({trees[750], lumberyards[750]}), .top_right({trees[751], lumberyards[751]}), .left(2'b0), .right({trees[801], lumberyards[801]}), .bottom_left(2'b0), .bottom({trees[850], lumberyards[850]}), .bottom_right({trees[851], lumberyards[851]}), .init(2'b00), .state({trees[800], lumberyards[800]}));
acre acre_16_1 (.clk(clk), .en(en), .top_left({trees[750], lumberyards[750]}), .top({trees[751], lumberyards[751]}), .top_right({trees[752], lumberyards[752]}), .left({trees[800], lumberyards[800]}), .right({trees[802], lumberyards[802]}), .bottom_left({trees[850], lumberyards[850]}), .bottom({trees[851], lumberyards[851]}), .bottom_right({trees[852], lumberyards[852]}), .init(2'b00), .state({trees[801], lumberyards[801]}));
acre acre_16_2 (.clk(clk), .en(en), .top_left({trees[751], lumberyards[751]}), .top({trees[752], lumberyards[752]}), .top_right({trees[753], lumberyards[753]}), .left({trees[801], lumberyards[801]}), .right({trees[803], lumberyards[803]}), .bottom_left({trees[851], lumberyards[851]}), .bottom({trees[852], lumberyards[852]}), .bottom_right({trees[853], lumberyards[853]}), .init(2'b00), .state({trees[802], lumberyards[802]}));
acre acre_16_3 (.clk(clk), .en(en), .top_left({trees[752], lumberyards[752]}), .top({trees[753], lumberyards[753]}), .top_right({trees[754], lumberyards[754]}), .left({trees[802], lumberyards[802]}), .right({trees[804], lumberyards[804]}), .bottom_left({trees[852], lumberyards[852]}), .bottom({trees[853], lumberyards[853]}), .bottom_right({trees[854], lumberyards[854]}), .init(2'b10), .state({trees[803], lumberyards[803]}));
acre acre_16_4 (.clk(clk), .en(en), .top_left({trees[753], lumberyards[753]}), .top({trees[754], lumberyards[754]}), .top_right({trees[755], lumberyards[755]}), .left({trees[803], lumberyards[803]}), .right({trees[805], lumberyards[805]}), .bottom_left({trees[853], lumberyards[853]}), .bottom({trees[854], lumberyards[854]}), .bottom_right({trees[855], lumberyards[855]}), .init(2'b00), .state({trees[804], lumberyards[804]}));
acre acre_16_5 (.clk(clk), .en(en), .top_left({trees[754], lumberyards[754]}), .top({trees[755], lumberyards[755]}), .top_right({trees[756], lumberyards[756]}), .left({trees[804], lumberyards[804]}), .right({trees[806], lumberyards[806]}), .bottom_left({trees[854], lumberyards[854]}), .bottom({trees[855], lumberyards[855]}), .bottom_right({trees[856], lumberyards[856]}), .init(2'b10), .state({trees[805], lumberyards[805]}));
acre acre_16_6 (.clk(clk), .en(en), .top_left({trees[755], lumberyards[755]}), .top({trees[756], lumberyards[756]}), .top_right({trees[757], lumberyards[757]}), .left({trees[805], lumberyards[805]}), .right({trees[807], lumberyards[807]}), .bottom_left({trees[855], lumberyards[855]}), .bottom({trees[856], lumberyards[856]}), .bottom_right({trees[857], lumberyards[857]}), .init(2'b01), .state({trees[806], lumberyards[806]}));
acre acre_16_7 (.clk(clk), .en(en), .top_left({trees[756], lumberyards[756]}), .top({trees[757], lumberyards[757]}), .top_right({trees[758], lumberyards[758]}), .left({trees[806], lumberyards[806]}), .right({trees[808], lumberyards[808]}), .bottom_left({trees[856], lumberyards[856]}), .bottom({trees[857], lumberyards[857]}), .bottom_right({trees[858], lumberyards[858]}), .init(2'b00), .state({trees[807], lumberyards[807]}));
acre acre_16_8 (.clk(clk), .en(en), .top_left({trees[757], lumberyards[757]}), .top({trees[758], lumberyards[758]}), .top_right({trees[759], lumberyards[759]}), .left({trees[807], lumberyards[807]}), .right({trees[809], lumberyards[809]}), .bottom_left({trees[857], lumberyards[857]}), .bottom({trees[858], lumberyards[858]}), .bottom_right({trees[859], lumberyards[859]}), .init(2'b00), .state({trees[808], lumberyards[808]}));
acre acre_16_9 (.clk(clk), .en(en), .top_left({trees[758], lumberyards[758]}), .top({trees[759], lumberyards[759]}), .top_right({trees[760], lumberyards[760]}), .left({trees[808], lumberyards[808]}), .right({trees[810], lumberyards[810]}), .bottom_left({trees[858], lumberyards[858]}), .bottom({trees[859], lumberyards[859]}), .bottom_right({trees[860], lumberyards[860]}), .init(2'b00), .state({trees[809], lumberyards[809]}));
acre acre_16_10 (.clk(clk), .en(en), .top_left({trees[759], lumberyards[759]}), .top({trees[760], lumberyards[760]}), .top_right({trees[761], lumberyards[761]}), .left({trees[809], lumberyards[809]}), .right({trees[811], lumberyards[811]}), .bottom_left({trees[859], lumberyards[859]}), .bottom({trees[860], lumberyards[860]}), .bottom_right({trees[861], lumberyards[861]}), .init(2'b00), .state({trees[810], lumberyards[810]}));
acre acre_16_11 (.clk(clk), .en(en), .top_left({trees[760], lumberyards[760]}), .top({trees[761], lumberyards[761]}), .top_right({trees[762], lumberyards[762]}), .left({trees[810], lumberyards[810]}), .right({trees[812], lumberyards[812]}), .bottom_left({trees[860], lumberyards[860]}), .bottom({trees[861], lumberyards[861]}), .bottom_right({trees[862], lumberyards[862]}), .init(2'b00), .state({trees[811], lumberyards[811]}));
acre acre_16_12 (.clk(clk), .en(en), .top_left({trees[761], lumberyards[761]}), .top({trees[762], lumberyards[762]}), .top_right({trees[763], lumberyards[763]}), .left({trees[811], lumberyards[811]}), .right({trees[813], lumberyards[813]}), .bottom_left({trees[861], lumberyards[861]}), .bottom({trees[862], lumberyards[862]}), .bottom_right({trees[863], lumberyards[863]}), .init(2'b00), .state({trees[812], lumberyards[812]}));
acre acre_16_13 (.clk(clk), .en(en), .top_left({trees[762], lumberyards[762]}), .top({trees[763], lumberyards[763]}), .top_right({trees[764], lumberyards[764]}), .left({trees[812], lumberyards[812]}), .right({trees[814], lumberyards[814]}), .bottom_left({trees[862], lumberyards[862]}), .bottom({trees[863], lumberyards[863]}), .bottom_right({trees[864], lumberyards[864]}), .init(2'b00), .state({trees[813], lumberyards[813]}));
acre acre_16_14 (.clk(clk), .en(en), .top_left({trees[763], lumberyards[763]}), .top({trees[764], lumberyards[764]}), .top_right({trees[765], lumberyards[765]}), .left({trees[813], lumberyards[813]}), .right({trees[815], lumberyards[815]}), .bottom_left({trees[863], lumberyards[863]}), .bottom({trees[864], lumberyards[864]}), .bottom_right({trees[865], lumberyards[865]}), .init(2'b00), .state({trees[814], lumberyards[814]}));
acre acre_16_15 (.clk(clk), .en(en), .top_left({trees[764], lumberyards[764]}), .top({trees[765], lumberyards[765]}), .top_right({trees[766], lumberyards[766]}), .left({trees[814], lumberyards[814]}), .right({trees[816], lumberyards[816]}), .bottom_left({trees[864], lumberyards[864]}), .bottom({trees[865], lumberyards[865]}), .bottom_right({trees[866], lumberyards[866]}), .init(2'b00), .state({trees[815], lumberyards[815]}));
acre acre_16_16 (.clk(clk), .en(en), .top_left({trees[765], lumberyards[765]}), .top({trees[766], lumberyards[766]}), .top_right({trees[767], lumberyards[767]}), .left({trees[815], lumberyards[815]}), .right({trees[817], lumberyards[817]}), .bottom_left({trees[865], lumberyards[865]}), .bottom({trees[866], lumberyards[866]}), .bottom_right({trees[867], lumberyards[867]}), .init(2'b00), .state({trees[816], lumberyards[816]}));
acre acre_16_17 (.clk(clk), .en(en), .top_left({trees[766], lumberyards[766]}), .top({trees[767], lumberyards[767]}), .top_right({trees[768], lumberyards[768]}), .left({trees[816], lumberyards[816]}), .right({trees[818], lumberyards[818]}), .bottom_left({trees[866], lumberyards[866]}), .bottom({trees[867], lumberyards[867]}), .bottom_right({trees[868], lumberyards[868]}), .init(2'b10), .state({trees[817], lumberyards[817]}));
acre acre_16_18 (.clk(clk), .en(en), .top_left({trees[767], lumberyards[767]}), .top({trees[768], lumberyards[768]}), .top_right({trees[769], lumberyards[769]}), .left({trees[817], lumberyards[817]}), .right({trees[819], lumberyards[819]}), .bottom_left({trees[867], lumberyards[867]}), .bottom({trees[868], lumberyards[868]}), .bottom_right({trees[869], lumberyards[869]}), .init(2'b00), .state({trees[818], lumberyards[818]}));
acre acre_16_19 (.clk(clk), .en(en), .top_left({trees[768], lumberyards[768]}), .top({trees[769], lumberyards[769]}), .top_right({trees[770], lumberyards[770]}), .left({trees[818], lumberyards[818]}), .right({trees[820], lumberyards[820]}), .bottom_left({trees[868], lumberyards[868]}), .bottom({trees[869], lumberyards[869]}), .bottom_right({trees[870], lumberyards[870]}), .init(2'b10), .state({trees[819], lumberyards[819]}));
acre acre_16_20 (.clk(clk), .en(en), .top_left({trees[769], lumberyards[769]}), .top({trees[770], lumberyards[770]}), .top_right({trees[771], lumberyards[771]}), .left({trees[819], lumberyards[819]}), .right({trees[821], lumberyards[821]}), .bottom_left({trees[869], lumberyards[869]}), .bottom({trees[870], lumberyards[870]}), .bottom_right({trees[871], lumberyards[871]}), .init(2'b00), .state({trees[820], lumberyards[820]}));
acre acre_16_21 (.clk(clk), .en(en), .top_left({trees[770], lumberyards[770]}), .top({trees[771], lumberyards[771]}), .top_right({trees[772], lumberyards[772]}), .left({trees[820], lumberyards[820]}), .right({trees[822], lumberyards[822]}), .bottom_left({trees[870], lumberyards[870]}), .bottom({trees[871], lumberyards[871]}), .bottom_right({trees[872], lumberyards[872]}), .init(2'b00), .state({trees[821], lumberyards[821]}));
acre acre_16_22 (.clk(clk), .en(en), .top_left({trees[771], lumberyards[771]}), .top({trees[772], lumberyards[772]}), .top_right({trees[773], lumberyards[773]}), .left({trees[821], lumberyards[821]}), .right({trees[823], lumberyards[823]}), .bottom_left({trees[871], lumberyards[871]}), .bottom({trees[872], lumberyards[872]}), .bottom_right({trees[873], lumberyards[873]}), .init(2'b10), .state({trees[822], lumberyards[822]}));
acre acre_16_23 (.clk(clk), .en(en), .top_left({trees[772], lumberyards[772]}), .top({trees[773], lumberyards[773]}), .top_right({trees[774], lumberyards[774]}), .left({trees[822], lumberyards[822]}), .right({trees[824], lumberyards[824]}), .bottom_left({trees[872], lumberyards[872]}), .bottom({trees[873], lumberyards[873]}), .bottom_right({trees[874], lumberyards[874]}), .init(2'b00), .state({trees[823], lumberyards[823]}));
acre acre_16_24 (.clk(clk), .en(en), .top_left({trees[773], lumberyards[773]}), .top({trees[774], lumberyards[774]}), .top_right({trees[775], lumberyards[775]}), .left({trees[823], lumberyards[823]}), .right({trees[825], lumberyards[825]}), .bottom_left({trees[873], lumberyards[873]}), .bottom({trees[874], lumberyards[874]}), .bottom_right({trees[875], lumberyards[875]}), .init(2'b00), .state({trees[824], lumberyards[824]}));
acre acre_16_25 (.clk(clk), .en(en), .top_left({trees[774], lumberyards[774]}), .top({trees[775], lumberyards[775]}), .top_right({trees[776], lumberyards[776]}), .left({trees[824], lumberyards[824]}), .right({trees[826], lumberyards[826]}), .bottom_left({trees[874], lumberyards[874]}), .bottom({trees[875], lumberyards[875]}), .bottom_right({trees[876], lumberyards[876]}), .init(2'b10), .state({trees[825], lumberyards[825]}));
acre acre_16_26 (.clk(clk), .en(en), .top_left({trees[775], lumberyards[775]}), .top({trees[776], lumberyards[776]}), .top_right({trees[777], lumberyards[777]}), .left({trees[825], lumberyards[825]}), .right({trees[827], lumberyards[827]}), .bottom_left({trees[875], lumberyards[875]}), .bottom({trees[876], lumberyards[876]}), .bottom_right({trees[877], lumberyards[877]}), .init(2'b00), .state({trees[826], lumberyards[826]}));
acre acre_16_27 (.clk(clk), .en(en), .top_left({trees[776], lumberyards[776]}), .top({trees[777], lumberyards[777]}), .top_right({trees[778], lumberyards[778]}), .left({trees[826], lumberyards[826]}), .right({trees[828], lumberyards[828]}), .bottom_left({trees[876], lumberyards[876]}), .bottom({trees[877], lumberyards[877]}), .bottom_right({trees[878], lumberyards[878]}), .init(2'b00), .state({trees[827], lumberyards[827]}));
acre acre_16_28 (.clk(clk), .en(en), .top_left({trees[777], lumberyards[777]}), .top({trees[778], lumberyards[778]}), .top_right({trees[779], lumberyards[779]}), .left({trees[827], lumberyards[827]}), .right({trees[829], lumberyards[829]}), .bottom_left({trees[877], lumberyards[877]}), .bottom({trees[878], lumberyards[878]}), .bottom_right({trees[879], lumberyards[879]}), .init(2'b00), .state({trees[828], lumberyards[828]}));
acre acre_16_29 (.clk(clk), .en(en), .top_left({trees[778], lumberyards[778]}), .top({trees[779], lumberyards[779]}), .top_right({trees[780], lumberyards[780]}), .left({trees[828], lumberyards[828]}), .right({trees[830], lumberyards[830]}), .bottom_left({trees[878], lumberyards[878]}), .bottom({trees[879], lumberyards[879]}), .bottom_right({trees[880], lumberyards[880]}), .init(2'b00), .state({trees[829], lumberyards[829]}));
acre acre_16_30 (.clk(clk), .en(en), .top_left({trees[779], lumberyards[779]}), .top({trees[780], lumberyards[780]}), .top_right({trees[781], lumberyards[781]}), .left({trees[829], lumberyards[829]}), .right({trees[831], lumberyards[831]}), .bottom_left({trees[879], lumberyards[879]}), .bottom({trees[880], lumberyards[880]}), .bottom_right({trees[881], lumberyards[881]}), .init(2'b00), .state({trees[830], lumberyards[830]}));
acre acre_16_31 (.clk(clk), .en(en), .top_left({trees[780], lumberyards[780]}), .top({trees[781], lumberyards[781]}), .top_right({trees[782], lumberyards[782]}), .left({trees[830], lumberyards[830]}), .right({trees[832], lumberyards[832]}), .bottom_left({trees[880], lumberyards[880]}), .bottom({trees[881], lumberyards[881]}), .bottom_right({trees[882], lumberyards[882]}), .init(2'b10), .state({trees[831], lumberyards[831]}));
acre acre_16_32 (.clk(clk), .en(en), .top_left({trees[781], lumberyards[781]}), .top({trees[782], lumberyards[782]}), .top_right({trees[783], lumberyards[783]}), .left({trees[831], lumberyards[831]}), .right({trees[833], lumberyards[833]}), .bottom_left({trees[881], lumberyards[881]}), .bottom({trees[882], lumberyards[882]}), .bottom_right({trees[883], lumberyards[883]}), .init(2'b00), .state({trees[832], lumberyards[832]}));
acre acre_16_33 (.clk(clk), .en(en), .top_left({trees[782], lumberyards[782]}), .top({trees[783], lumberyards[783]}), .top_right({trees[784], lumberyards[784]}), .left({trees[832], lumberyards[832]}), .right({trees[834], lumberyards[834]}), .bottom_left({trees[882], lumberyards[882]}), .bottom({trees[883], lumberyards[883]}), .bottom_right({trees[884], lumberyards[884]}), .init(2'b01), .state({trees[833], lumberyards[833]}));
acre acre_16_34 (.clk(clk), .en(en), .top_left({trees[783], lumberyards[783]}), .top({trees[784], lumberyards[784]}), .top_right({trees[785], lumberyards[785]}), .left({trees[833], lumberyards[833]}), .right({trees[835], lumberyards[835]}), .bottom_left({trees[883], lumberyards[883]}), .bottom({trees[884], lumberyards[884]}), .bottom_right({trees[885], lumberyards[885]}), .init(2'b10), .state({trees[834], lumberyards[834]}));
acre acre_16_35 (.clk(clk), .en(en), .top_left({trees[784], lumberyards[784]}), .top({trees[785], lumberyards[785]}), .top_right({trees[786], lumberyards[786]}), .left({trees[834], lumberyards[834]}), .right({trees[836], lumberyards[836]}), .bottom_left({trees[884], lumberyards[884]}), .bottom({trees[885], lumberyards[885]}), .bottom_right({trees[886], lumberyards[886]}), .init(2'b00), .state({trees[835], lumberyards[835]}));
acre acre_16_36 (.clk(clk), .en(en), .top_left({trees[785], lumberyards[785]}), .top({trees[786], lumberyards[786]}), .top_right({trees[787], lumberyards[787]}), .left({trees[835], lumberyards[835]}), .right({trees[837], lumberyards[837]}), .bottom_left({trees[885], lumberyards[885]}), .bottom({trees[886], lumberyards[886]}), .bottom_right({trees[887], lumberyards[887]}), .init(2'b00), .state({trees[836], lumberyards[836]}));
acre acre_16_37 (.clk(clk), .en(en), .top_left({trees[786], lumberyards[786]}), .top({trees[787], lumberyards[787]}), .top_right({trees[788], lumberyards[788]}), .left({trees[836], lumberyards[836]}), .right({trees[838], lumberyards[838]}), .bottom_left({trees[886], lumberyards[886]}), .bottom({trees[887], lumberyards[887]}), .bottom_right({trees[888], lumberyards[888]}), .init(2'b01), .state({trees[837], lumberyards[837]}));
acre acre_16_38 (.clk(clk), .en(en), .top_left({trees[787], lumberyards[787]}), .top({trees[788], lumberyards[788]}), .top_right({trees[789], lumberyards[789]}), .left({trees[837], lumberyards[837]}), .right({trees[839], lumberyards[839]}), .bottom_left({trees[887], lumberyards[887]}), .bottom({trees[888], lumberyards[888]}), .bottom_right({trees[889], lumberyards[889]}), .init(2'b10), .state({trees[838], lumberyards[838]}));
acre acre_16_39 (.clk(clk), .en(en), .top_left({trees[788], lumberyards[788]}), .top({trees[789], lumberyards[789]}), .top_right({trees[790], lumberyards[790]}), .left({trees[838], lumberyards[838]}), .right({trees[840], lumberyards[840]}), .bottom_left({trees[888], lumberyards[888]}), .bottom({trees[889], lumberyards[889]}), .bottom_right({trees[890], lumberyards[890]}), .init(2'b00), .state({trees[839], lumberyards[839]}));
acre acre_16_40 (.clk(clk), .en(en), .top_left({trees[789], lumberyards[789]}), .top({trees[790], lumberyards[790]}), .top_right({trees[791], lumberyards[791]}), .left({trees[839], lumberyards[839]}), .right({trees[841], lumberyards[841]}), .bottom_left({trees[889], lumberyards[889]}), .bottom({trees[890], lumberyards[890]}), .bottom_right({trees[891], lumberyards[891]}), .init(2'b00), .state({trees[840], lumberyards[840]}));
acre acre_16_41 (.clk(clk), .en(en), .top_left({trees[790], lumberyards[790]}), .top({trees[791], lumberyards[791]}), .top_right({trees[792], lumberyards[792]}), .left({trees[840], lumberyards[840]}), .right({trees[842], lumberyards[842]}), .bottom_left({trees[890], lumberyards[890]}), .bottom({trees[891], lumberyards[891]}), .bottom_right({trees[892], lumberyards[892]}), .init(2'b00), .state({trees[841], lumberyards[841]}));
acre acre_16_42 (.clk(clk), .en(en), .top_left({trees[791], lumberyards[791]}), .top({trees[792], lumberyards[792]}), .top_right({trees[793], lumberyards[793]}), .left({trees[841], lumberyards[841]}), .right({trees[843], lumberyards[843]}), .bottom_left({trees[891], lumberyards[891]}), .bottom({trees[892], lumberyards[892]}), .bottom_right({trees[893], lumberyards[893]}), .init(2'b10), .state({trees[842], lumberyards[842]}));
acre acre_16_43 (.clk(clk), .en(en), .top_left({trees[792], lumberyards[792]}), .top({trees[793], lumberyards[793]}), .top_right({trees[794], lumberyards[794]}), .left({trees[842], lumberyards[842]}), .right({trees[844], lumberyards[844]}), .bottom_left({trees[892], lumberyards[892]}), .bottom({trees[893], lumberyards[893]}), .bottom_right({trees[894], lumberyards[894]}), .init(2'b00), .state({trees[843], lumberyards[843]}));
acre acre_16_44 (.clk(clk), .en(en), .top_left({trees[793], lumberyards[793]}), .top({trees[794], lumberyards[794]}), .top_right({trees[795], lumberyards[795]}), .left({trees[843], lumberyards[843]}), .right({trees[845], lumberyards[845]}), .bottom_left({trees[893], lumberyards[893]}), .bottom({trees[894], lumberyards[894]}), .bottom_right({trees[895], lumberyards[895]}), .init(2'b00), .state({trees[844], lumberyards[844]}));
acre acre_16_45 (.clk(clk), .en(en), .top_left({trees[794], lumberyards[794]}), .top({trees[795], lumberyards[795]}), .top_right({trees[796], lumberyards[796]}), .left({trees[844], lumberyards[844]}), .right({trees[846], lumberyards[846]}), .bottom_left({trees[894], lumberyards[894]}), .bottom({trees[895], lumberyards[895]}), .bottom_right({trees[896], lumberyards[896]}), .init(2'b00), .state({trees[845], lumberyards[845]}));
acre acre_16_46 (.clk(clk), .en(en), .top_left({trees[795], lumberyards[795]}), .top({trees[796], lumberyards[796]}), .top_right({trees[797], lumberyards[797]}), .left({trees[845], lumberyards[845]}), .right({trees[847], lumberyards[847]}), .bottom_left({trees[895], lumberyards[895]}), .bottom({trees[896], lumberyards[896]}), .bottom_right({trees[897], lumberyards[897]}), .init(2'b10), .state({trees[846], lumberyards[846]}));
acre acre_16_47 (.clk(clk), .en(en), .top_left({trees[796], lumberyards[796]}), .top({trees[797], lumberyards[797]}), .top_right({trees[798], lumberyards[798]}), .left({trees[846], lumberyards[846]}), .right({trees[848], lumberyards[848]}), .bottom_left({trees[896], lumberyards[896]}), .bottom({trees[897], lumberyards[897]}), .bottom_right({trees[898], lumberyards[898]}), .init(2'b00), .state({trees[847], lumberyards[847]}));
acre acre_16_48 (.clk(clk), .en(en), .top_left({trees[797], lumberyards[797]}), .top({trees[798], lumberyards[798]}), .top_right({trees[799], lumberyards[799]}), .left({trees[847], lumberyards[847]}), .right({trees[849], lumberyards[849]}), .bottom_left({trees[897], lumberyards[897]}), .bottom({trees[898], lumberyards[898]}), .bottom_right({trees[899], lumberyards[899]}), .init(2'b00), .state({trees[848], lumberyards[848]}));
acre acre_16_49 (.clk(clk), .en(en), .top_left({trees[798], lumberyards[798]}), .top({trees[799], lumberyards[799]}), .top_right(2'b0), .left({trees[848], lumberyards[848]}), .right(2'b0), .bottom_left({trees[898], lumberyards[898]}), .bottom({trees[899], lumberyards[899]}), .bottom_right(2'b0), .init(2'b01), .state({trees[849], lumberyards[849]}));
acre acre_17_0 (.clk(clk), .en(en), .top_left(2'b0), .top({trees[800], lumberyards[800]}), .top_right({trees[801], lumberyards[801]}), .left(2'b0), .right({trees[851], lumberyards[851]}), .bottom_left(2'b0), .bottom({trees[900], lumberyards[900]}), .bottom_right({trees[901], lumberyards[901]}), .init(2'b00), .state({trees[850], lumberyards[850]}));
acre acre_17_1 (.clk(clk), .en(en), .top_left({trees[800], lumberyards[800]}), .top({trees[801], lumberyards[801]}), .top_right({trees[802], lumberyards[802]}), .left({trees[850], lumberyards[850]}), .right({trees[852], lumberyards[852]}), .bottom_left({trees[900], lumberyards[900]}), .bottom({trees[901], lumberyards[901]}), .bottom_right({trees[902], lumberyards[902]}), .init(2'b00), .state({trees[851], lumberyards[851]}));
acre acre_17_2 (.clk(clk), .en(en), .top_left({trees[801], lumberyards[801]}), .top({trees[802], lumberyards[802]}), .top_right({trees[803], lumberyards[803]}), .left({trees[851], lumberyards[851]}), .right({trees[853], lumberyards[853]}), .bottom_left({trees[901], lumberyards[901]}), .bottom({trees[902], lumberyards[902]}), .bottom_right({trees[903], lumberyards[903]}), .init(2'b01), .state({trees[852], lumberyards[852]}));
acre acre_17_3 (.clk(clk), .en(en), .top_left({trees[802], lumberyards[802]}), .top({trees[803], lumberyards[803]}), .top_right({trees[804], lumberyards[804]}), .left({trees[852], lumberyards[852]}), .right({trees[854], lumberyards[854]}), .bottom_left({trees[902], lumberyards[902]}), .bottom({trees[903], lumberyards[903]}), .bottom_right({trees[904], lumberyards[904]}), .init(2'b00), .state({trees[853], lumberyards[853]}));
acre acre_17_4 (.clk(clk), .en(en), .top_left({trees[803], lumberyards[803]}), .top({trees[804], lumberyards[804]}), .top_right({trees[805], lumberyards[805]}), .left({trees[853], lumberyards[853]}), .right({trees[855], lumberyards[855]}), .bottom_left({trees[903], lumberyards[903]}), .bottom({trees[904], lumberyards[904]}), .bottom_right({trees[905], lumberyards[905]}), .init(2'b00), .state({trees[854], lumberyards[854]}));
acre acre_17_5 (.clk(clk), .en(en), .top_left({trees[804], lumberyards[804]}), .top({trees[805], lumberyards[805]}), .top_right({trees[806], lumberyards[806]}), .left({trees[854], lumberyards[854]}), .right({trees[856], lumberyards[856]}), .bottom_left({trees[904], lumberyards[904]}), .bottom({trees[905], lumberyards[905]}), .bottom_right({trees[906], lumberyards[906]}), .init(2'b00), .state({trees[855], lumberyards[855]}));
acre acre_17_6 (.clk(clk), .en(en), .top_left({trees[805], lumberyards[805]}), .top({trees[806], lumberyards[806]}), .top_right({trees[807], lumberyards[807]}), .left({trees[855], lumberyards[855]}), .right({trees[857], lumberyards[857]}), .bottom_left({trees[905], lumberyards[905]}), .bottom({trees[906], lumberyards[906]}), .bottom_right({trees[907], lumberyards[907]}), .init(2'b10), .state({trees[856], lumberyards[856]}));
acre acre_17_7 (.clk(clk), .en(en), .top_left({trees[806], lumberyards[806]}), .top({trees[807], lumberyards[807]}), .top_right({trees[808], lumberyards[808]}), .left({trees[856], lumberyards[856]}), .right({trees[858], lumberyards[858]}), .bottom_left({trees[906], lumberyards[906]}), .bottom({trees[907], lumberyards[907]}), .bottom_right({trees[908], lumberyards[908]}), .init(2'b00), .state({trees[857], lumberyards[857]}));
acre acre_17_8 (.clk(clk), .en(en), .top_left({trees[807], lumberyards[807]}), .top({trees[808], lumberyards[808]}), .top_right({trees[809], lumberyards[809]}), .left({trees[857], lumberyards[857]}), .right({trees[859], lumberyards[859]}), .bottom_left({trees[907], lumberyards[907]}), .bottom({trees[908], lumberyards[908]}), .bottom_right({trees[909], lumberyards[909]}), .init(2'b00), .state({trees[858], lumberyards[858]}));
acre acre_17_9 (.clk(clk), .en(en), .top_left({trees[808], lumberyards[808]}), .top({trees[809], lumberyards[809]}), .top_right({trees[810], lumberyards[810]}), .left({trees[858], lumberyards[858]}), .right({trees[860], lumberyards[860]}), .bottom_left({trees[908], lumberyards[908]}), .bottom({trees[909], lumberyards[909]}), .bottom_right({trees[910], lumberyards[910]}), .init(2'b00), .state({trees[859], lumberyards[859]}));
acre acre_17_10 (.clk(clk), .en(en), .top_left({trees[809], lumberyards[809]}), .top({trees[810], lumberyards[810]}), .top_right({trees[811], lumberyards[811]}), .left({trees[859], lumberyards[859]}), .right({trees[861], lumberyards[861]}), .bottom_left({trees[909], lumberyards[909]}), .bottom({trees[910], lumberyards[910]}), .bottom_right({trees[911], lumberyards[911]}), .init(2'b01), .state({trees[860], lumberyards[860]}));
acre acre_17_11 (.clk(clk), .en(en), .top_left({trees[810], lumberyards[810]}), .top({trees[811], lumberyards[811]}), .top_right({trees[812], lumberyards[812]}), .left({trees[860], lumberyards[860]}), .right({trees[862], lumberyards[862]}), .bottom_left({trees[910], lumberyards[910]}), .bottom({trees[911], lumberyards[911]}), .bottom_right({trees[912], lumberyards[912]}), .init(2'b00), .state({trees[861], lumberyards[861]}));
acre acre_17_12 (.clk(clk), .en(en), .top_left({trees[811], lumberyards[811]}), .top({trees[812], lumberyards[812]}), .top_right({trees[813], lumberyards[813]}), .left({trees[861], lumberyards[861]}), .right({trees[863], lumberyards[863]}), .bottom_left({trees[911], lumberyards[911]}), .bottom({trees[912], lumberyards[912]}), .bottom_right({trees[913], lumberyards[913]}), .init(2'b01), .state({trees[862], lumberyards[862]}));
acre acre_17_13 (.clk(clk), .en(en), .top_left({trees[812], lumberyards[812]}), .top({trees[813], lumberyards[813]}), .top_right({trees[814], lumberyards[814]}), .left({trees[862], lumberyards[862]}), .right({trees[864], lumberyards[864]}), .bottom_left({trees[912], lumberyards[912]}), .bottom({trees[913], lumberyards[913]}), .bottom_right({trees[914], lumberyards[914]}), .init(2'b10), .state({trees[863], lumberyards[863]}));
acre acre_17_14 (.clk(clk), .en(en), .top_left({trees[813], lumberyards[813]}), .top({trees[814], lumberyards[814]}), .top_right({trees[815], lumberyards[815]}), .left({trees[863], lumberyards[863]}), .right({trees[865], lumberyards[865]}), .bottom_left({trees[913], lumberyards[913]}), .bottom({trees[914], lumberyards[914]}), .bottom_right({trees[915], lumberyards[915]}), .init(2'b10), .state({trees[864], lumberyards[864]}));
acre acre_17_15 (.clk(clk), .en(en), .top_left({trees[814], lumberyards[814]}), .top({trees[815], lumberyards[815]}), .top_right({trees[816], lumberyards[816]}), .left({trees[864], lumberyards[864]}), .right({trees[866], lumberyards[866]}), .bottom_left({trees[914], lumberyards[914]}), .bottom({trees[915], lumberyards[915]}), .bottom_right({trees[916], lumberyards[916]}), .init(2'b00), .state({trees[865], lumberyards[865]}));
acre acre_17_16 (.clk(clk), .en(en), .top_left({trees[815], lumberyards[815]}), .top({trees[816], lumberyards[816]}), .top_right({trees[817], lumberyards[817]}), .left({trees[865], lumberyards[865]}), .right({trees[867], lumberyards[867]}), .bottom_left({trees[915], lumberyards[915]}), .bottom({trees[916], lumberyards[916]}), .bottom_right({trees[917], lumberyards[917]}), .init(2'b00), .state({trees[866], lumberyards[866]}));
acre acre_17_17 (.clk(clk), .en(en), .top_left({trees[816], lumberyards[816]}), .top({trees[817], lumberyards[817]}), .top_right({trees[818], lumberyards[818]}), .left({trees[866], lumberyards[866]}), .right({trees[868], lumberyards[868]}), .bottom_left({trees[916], lumberyards[916]}), .bottom({trees[917], lumberyards[917]}), .bottom_right({trees[918], lumberyards[918]}), .init(2'b00), .state({trees[867], lumberyards[867]}));
acre acre_17_18 (.clk(clk), .en(en), .top_left({trees[817], lumberyards[817]}), .top({trees[818], lumberyards[818]}), .top_right({trees[819], lumberyards[819]}), .left({trees[867], lumberyards[867]}), .right({trees[869], lumberyards[869]}), .bottom_left({trees[917], lumberyards[917]}), .bottom({trees[918], lumberyards[918]}), .bottom_right({trees[919], lumberyards[919]}), .init(2'b01), .state({trees[868], lumberyards[868]}));
acre acre_17_19 (.clk(clk), .en(en), .top_left({trees[818], lumberyards[818]}), .top({trees[819], lumberyards[819]}), .top_right({trees[820], lumberyards[820]}), .left({trees[868], lumberyards[868]}), .right({trees[870], lumberyards[870]}), .bottom_left({trees[918], lumberyards[918]}), .bottom({trees[919], lumberyards[919]}), .bottom_right({trees[920], lumberyards[920]}), .init(2'b00), .state({trees[869], lumberyards[869]}));
acre acre_17_20 (.clk(clk), .en(en), .top_left({trees[819], lumberyards[819]}), .top({trees[820], lumberyards[820]}), .top_right({trees[821], lumberyards[821]}), .left({trees[869], lumberyards[869]}), .right({trees[871], lumberyards[871]}), .bottom_left({trees[919], lumberyards[919]}), .bottom({trees[920], lumberyards[920]}), .bottom_right({trees[921], lumberyards[921]}), .init(2'b00), .state({trees[870], lumberyards[870]}));
acre acre_17_21 (.clk(clk), .en(en), .top_left({trees[820], lumberyards[820]}), .top({trees[821], lumberyards[821]}), .top_right({trees[822], lumberyards[822]}), .left({trees[870], lumberyards[870]}), .right({trees[872], lumberyards[872]}), .bottom_left({trees[920], lumberyards[920]}), .bottom({trees[921], lumberyards[921]}), .bottom_right({trees[922], lumberyards[922]}), .init(2'b10), .state({trees[871], lumberyards[871]}));
acre acre_17_22 (.clk(clk), .en(en), .top_left({trees[821], lumberyards[821]}), .top({trees[822], lumberyards[822]}), .top_right({trees[823], lumberyards[823]}), .left({trees[871], lumberyards[871]}), .right({trees[873], lumberyards[873]}), .bottom_left({trees[921], lumberyards[921]}), .bottom({trees[922], lumberyards[922]}), .bottom_right({trees[923], lumberyards[923]}), .init(2'b00), .state({trees[872], lumberyards[872]}));
acre acre_17_23 (.clk(clk), .en(en), .top_left({trees[822], lumberyards[822]}), .top({trees[823], lumberyards[823]}), .top_right({trees[824], lumberyards[824]}), .left({trees[872], lumberyards[872]}), .right({trees[874], lumberyards[874]}), .bottom_left({trees[922], lumberyards[922]}), .bottom({trees[923], lumberyards[923]}), .bottom_right({trees[924], lumberyards[924]}), .init(2'b00), .state({trees[873], lumberyards[873]}));
acre acre_17_24 (.clk(clk), .en(en), .top_left({trees[823], lumberyards[823]}), .top({trees[824], lumberyards[824]}), .top_right({trees[825], lumberyards[825]}), .left({trees[873], lumberyards[873]}), .right({trees[875], lumberyards[875]}), .bottom_left({trees[923], lumberyards[923]}), .bottom({trees[924], lumberyards[924]}), .bottom_right({trees[925], lumberyards[925]}), .init(2'b01), .state({trees[874], lumberyards[874]}));
acre acre_17_25 (.clk(clk), .en(en), .top_left({trees[824], lumberyards[824]}), .top({trees[825], lumberyards[825]}), .top_right({trees[826], lumberyards[826]}), .left({trees[874], lumberyards[874]}), .right({trees[876], lumberyards[876]}), .bottom_left({trees[924], lumberyards[924]}), .bottom({trees[925], lumberyards[925]}), .bottom_right({trees[926], lumberyards[926]}), .init(2'b10), .state({trees[875], lumberyards[875]}));
acre acre_17_26 (.clk(clk), .en(en), .top_left({trees[825], lumberyards[825]}), .top({trees[826], lumberyards[826]}), .top_right({trees[827], lumberyards[827]}), .left({trees[875], lumberyards[875]}), .right({trees[877], lumberyards[877]}), .bottom_left({trees[925], lumberyards[925]}), .bottom({trees[926], lumberyards[926]}), .bottom_right({trees[927], lumberyards[927]}), .init(2'b01), .state({trees[876], lumberyards[876]}));
acre acre_17_27 (.clk(clk), .en(en), .top_left({trees[826], lumberyards[826]}), .top({trees[827], lumberyards[827]}), .top_right({trees[828], lumberyards[828]}), .left({trees[876], lumberyards[876]}), .right({trees[878], lumberyards[878]}), .bottom_left({trees[926], lumberyards[926]}), .bottom({trees[927], lumberyards[927]}), .bottom_right({trees[928], lumberyards[928]}), .init(2'b00), .state({trees[877], lumberyards[877]}));
acre acre_17_28 (.clk(clk), .en(en), .top_left({trees[827], lumberyards[827]}), .top({trees[828], lumberyards[828]}), .top_right({trees[829], lumberyards[829]}), .left({trees[877], lumberyards[877]}), .right({trees[879], lumberyards[879]}), .bottom_left({trees[927], lumberyards[927]}), .bottom({trees[928], lumberyards[928]}), .bottom_right({trees[929], lumberyards[929]}), .init(2'b00), .state({trees[878], lumberyards[878]}));
acre acre_17_29 (.clk(clk), .en(en), .top_left({trees[828], lumberyards[828]}), .top({trees[829], lumberyards[829]}), .top_right({trees[830], lumberyards[830]}), .left({trees[878], lumberyards[878]}), .right({trees[880], lumberyards[880]}), .bottom_left({trees[928], lumberyards[928]}), .bottom({trees[929], lumberyards[929]}), .bottom_right({trees[930], lumberyards[930]}), .init(2'b00), .state({trees[879], lumberyards[879]}));
acre acre_17_30 (.clk(clk), .en(en), .top_left({trees[829], lumberyards[829]}), .top({trees[830], lumberyards[830]}), .top_right({trees[831], lumberyards[831]}), .left({trees[879], lumberyards[879]}), .right({trees[881], lumberyards[881]}), .bottom_left({trees[929], lumberyards[929]}), .bottom({trees[930], lumberyards[930]}), .bottom_right({trees[931], lumberyards[931]}), .init(2'b00), .state({trees[880], lumberyards[880]}));
acre acre_17_31 (.clk(clk), .en(en), .top_left({trees[830], lumberyards[830]}), .top({trees[831], lumberyards[831]}), .top_right({trees[832], lumberyards[832]}), .left({trees[880], lumberyards[880]}), .right({trees[882], lumberyards[882]}), .bottom_left({trees[930], lumberyards[930]}), .bottom({trees[931], lumberyards[931]}), .bottom_right({trees[932], lumberyards[932]}), .init(2'b01), .state({trees[881], lumberyards[881]}));
acre acre_17_32 (.clk(clk), .en(en), .top_left({trees[831], lumberyards[831]}), .top({trees[832], lumberyards[832]}), .top_right({trees[833], lumberyards[833]}), .left({trees[881], lumberyards[881]}), .right({trees[883], lumberyards[883]}), .bottom_left({trees[931], lumberyards[931]}), .bottom({trees[932], lumberyards[932]}), .bottom_right({trees[933], lumberyards[933]}), .init(2'b01), .state({trees[882], lumberyards[882]}));
acre acre_17_33 (.clk(clk), .en(en), .top_left({trees[832], lumberyards[832]}), .top({trees[833], lumberyards[833]}), .top_right({trees[834], lumberyards[834]}), .left({trees[882], lumberyards[882]}), .right({trees[884], lumberyards[884]}), .bottom_left({trees[932], lumberyards[932]}), .bottom({trees[933], lumberyards[933]}), .bottom_right({trees[934], lumberyards[934]}), .init(2'b00), .state({trees[883], lumberyards[883]}));
acre acre_17_34 (.clk(clk), .en(en), .top_left({trees[833], lumberyards[833]}), .top({trees[834], lumberyards[834]}), .top_right({trees[835], lumberyards[835]}), .left({trees[883], lumberyards[883]}), .right({trees[885], lumberyards[885]}), .bottom_left({trees[933], lumberyards[933]}), .bottom({trees[934], lumberyards[934]}), .bottom_right({trees[935], lumberyards[935]}), .init(2'b00), .state({trees[884], lumberyards[884]}));
acre acre_17_35 (.clk(clk), .en(en), .top_left({trees[834], lumberyards[834]}), .top({trees[835], lumberyards[835]}), .top_right({trees[836], lumberyards[836]}), .left({trees[884], lumberyards[884]}), .right({trees[886], lumberyards[886]}), .bottom_left({trees[934], lumberyards[934]}), .bottom({trees[935], lumberyards[935]}), .bottom_right({trees[936], lumberyards[936]}), .init(2'b01), .state({trees[885], lumberyards[885]}));
acre acre_17_36 (.clk(clk), .en(en), .top_left({trees[835], lumberyards[835]}), .top({trees[836], lumberyards[836]}), .top_right({trees[837], lumberyards[837]}), .left({trees[885], lumberyards[885]}), .right({trees[887], lumberyards[887]}), .bottom_left({trees[935], lumberyards[935]}), .bottom({trees[936], lumberyards[936]}), .bottom_right({trees[937], lumberyards[937]}), .init(2'b00), .state({trees[886], lumberyards[886]}));
acre acre_17_37 (.clk(clk), .en(en), .top_left({trees[836], lumberyards[836]}), .top({trees[837], lumberyards[837]}), .top_right({trees[838], lumberyards[838]}), .left({trees[886], lumberyards[886]}), .right({trees[888], lumberyards[888]}), .bottom_left({trees[936], lumberyards[936]}), .bottom({trees[937], lumberyards[937]}), .bottom_right({trees[938], lumberyards[938]}), .init(2'b00), .state({trees[887], lumberyards[887]}));
acre acre_17_38 (.clk(clk), .en(en), .top_left({trees[837], lumberyards[837]}), .top({trees[838], lumberyards[838]}), .top_right({trees[839], lumberyards[839]}), .left({trees[887], lumberyards[887]}), .right({trees[889], lumberyards[889]}), .bottom_left({trees[937], lumberyards[937]}), .bottom({trees[938], lumberyards[938]}), .bottom_right({trees[939], lumberyards[939]}), .init(2'b00), .state({trees[888], lumberyards[888]}));
acre acre_17_39 (.clk(clk), .en(en), .top_left({trees[838], lumberyards[838]}), .top({trees[839], lumberyards[839]}), .top_right({trees[840], lumberyards[840]}), .left({trees[888], lumberyards[888]}), .right({trees[890], lumberyards[890]}), .bottom_left({trees[938], lumberyards[938]}), .bottom({trees[939], lumberyards[939]}), .bottom_right({trees[940], lumberyards[940]}), .init(2'b00), .state({trees[889], lumberyards[889]}));
acre acre_17_40 (.clk(clk), .en(en), .top_left({trees[839], lumberyards[839]}), .top({trees[840], lumberyards[840]}), .top_right({trees[841], lumberyards[841]}), .left({trees[889], lumberyards[889]}), .right({trees[891], lumberyards[891]}), .bottom_left({trees[939], lumberyards[939]}), .bottom({trees[940], lumberyards[940]}), .bottom_right({trees[941], lumberyards[941]}), .init(2'b00), .state({trees[890], lumberyards[890]}));
acre acre_17_41 (.clk(clk), .en(en), .top_left({trees[840], lumberyards[840]}), .top({trees[841], lumberyards[841]}), .top_right({trees[842], lumberyards[842]}), .left({trees[890], lumberyards[890]}), .right({trees[892], lumberyards[892]}), .bottom_left({trees[940], lumberyards[940]}), .bottom({trees[941], lumberyards[941]}), .bottom_right({trees[942], lumberyards[942]}), .init(2'b00), .state({trees[891], lumberyards[891]}));
acre acre_17_42 (.clk(clk), .en(en), .top_left({trees[841], lumberyards[841]}), .top({trees[842], lumberyards[842]}), .top_right({trees[843], lumberyards[843]}), .left({trees[891], lumberyards[891]}), .right({trees[893], lumberyards[893]}), .bottom_left({trees[941], lumberyards[941]}), .bottom({trees[942], lumberyards[942]}), .bottom_right({trees[943], lumberyards[943]}), .init(2'b01), .state({trees[892], lumberyards[892]}));
acre acre_17_43 (.clk(clk), .en(en), .top_left({trees[842], lumberyards[842]}), .top({trees[843], lumberyards[843]}), .top_right({trees[844], lumberyards[844]}), .left({trees[892], lumberyards[892]}), .right({trees[894], lumberyards[894]}), .bottom_left({trees[942], lumberyards[942]}), .bottom({trees[943], lumberyards[943]}), .bottom_right({trees[944], lumberyards[944]}), .init(2'b01), .state({trees[893], lumberyards[893]}));
acre acre_17_44 (.clk(clk), .en(en), .top_left({trees[843], lumberyards[843]}), .top({trees[844], lumberyards[844]}), .top_right({trees[845], lumberyards[845]}), .left({trees[893], lumberyards[893]}), .right({trees[895], lumberyards[895]}), .bottom_left({trees[943], lumberyards[943]}), .bottom({trees[944], lumberyards[944]}), .bottom_right({trees[945], lumberyards[945]}), .init(2'b01), .state({trees[894], lumberyards[894]}));
acre acre_17_45 (.clk(clk), .en(en), .top_left({trees[844], lumberyards[844]}), .top({trees[845], lumberyards[845]}), .top_right({trees[846], lumberyards[846]}), .left({trees[894], lumberyards[894]}), .right({trees[896], lumberyards[896]}), .bottom_left({trees[944], lumberyards[944]}), .bottom({trees[945], lumberyards[945]}), .bottom_right({trees[946], lumberyards[946]}), .init(2'b01), .state({trees[895], lumberyards[895]}));
acre acre_17_46 (.clk(clk), .en(en), .top_left({trees[845], lumberyards[845]}), .top({trees[846], lumberyards[846]}), .top_right({trees[847], lumberyards[847]}), .left({trees[895], lumberyards[895]}), .right({trees[897], lumberyards[897]}), .bottom_left({trees[945], lumberyards[945]}), .bottom({trees[946], lumberyards[946]}), .bottom_right({trees[947], lumberyards[947]}), .init(2'b00), .state({trees[896], lumberyards[896]}));
acre acre_17_47 (.clk(clk), .en(en), .top_left({trees[846], lumberyards[846]}), .top({trees[847], lumberyards[847]}), .top_right({trees[848], lumberyards[848]}), .left({trees[896], lumberyards[896]}), .right({trees[898], lumberyards[898]}), .bottom_left({trees[946], lumberyards[946]}), .bottom({trees[947], lumberyards[947]}), .bottom_right({trees[948], lumberyards[948]}), .init(2'b00), .state({trees[897], lumberyards[897]}));
acre acre_17_48 (.clk(clk), .en(en), .top_left({trees[847], lumberyards[847]}), .top({trees[848], lumberyards[848]}), .top_right({trees[849], lumberyards[849]}), .left({trees[897], lumberyards[897]}), .right({trees[899], lumberyards[899]}), .bottom_left({trees[947], lumberyards[947]}), .bottom({trees[948], lumberyards[948]}), .bottom_right({trees[949], lumberyards[949]}), .init(2'b10), .state({trees[898], lumberyards[898]}));
acre acre_17_49 (.clk(clk), .en(en), .top_left({trees[848], lumberyards[848]}), .top({trees[849], lumberyards[849]}), .top_right(2'b0), .left({trees[898], lumberyards[898]}), .right(2'b0), .bottom_left({trees[948], lumberyards[948]}), .bottom({trees[949], lumberyards[949]}), .bottom_right(2'b0), .init(2'b00), .state({trees[899], lumberyards[899]}));
acre acre_18_0 (.clk(clk), .en(en), .top_left(2'b0), .top({trees[850], lumberyards[850]}), .top_right({trees[851], lumberyards[851]}), .left(2'b0), .right({trees[901], lumberyards[901]}), .bottom_left(2'b0), .bottom({trees[950], lumberyards[950]}), .bottom_right({trees[951], lumberyards[951]}), .init(2'b00), .state({trees[900], lumberyards[900]}));
acre acre_18_1 (.clk(clk), .en(en), .top_left({trees[850], lumberyards[850]}), .top({trees[851], lumberyards[851]}), .top_right({trees[852], lumberyards[852]}), .left({trees[900], lumberyards[900]}), .right({trees[902], lumberyards[902]}), .bottom_left({trees[950], lumberyards[950]}), .bottom({trees[951], lumberyards[951]}), .bottom_right({trees[952], lumberyards[952]}), .init(2'b00), .state({trees[901], lumberyards[901]}));
acre acre_18_2 (.clk(clk), .en(en), .top_left({trees[851], lumberyards[851]}), .top({trees[852], lumberyards[852]}), .top_right({trees[853], lumberyards[853]}), .left({trees[901], lumberyards[901]}), .right({trees[903], lumberyards[903]}), .bottom_left({trees[951], lumberyards[951]}), .bottom({trees[952], lumberyards[952]}), .bottom_right({trees[953], lumberyards[953]}), .init(2'b00), .state({trees[902], lumberyards[902]}));
acre acre_18_3 (.clk(clk), .en(en), .top_left({trees[852], lumberyards[852]}), .top({trees[853], lumberyards[853]}), .top_right({trees[854], lumberyards[854]}), .left({trees[902], lumberyards[902]}), .right({trees[904], lumberyards[904]}), .bottom_left({trees[952], lumberyards[952]}), .bottom({trees[953], lumberyards[953]}), .bottom_right({trees[954], lumberyards[954]}), .init(2'b00), .state({trees[903], lumberyards[903]}));
acre acre_18_4 (.clk(clk), .en(en), .top_left({trees[853], lumberyards[853]}), .top({trees[854], lumberyards[854]}), .top_right({trees[855], lumberyards[855]}), .left({trees[903], lumberyards[903]}), .right({trees[905], lumberyards[905]}), .bottom_left({trees[953], lumberyards[953]}), .bottom({trees[954], lumberyards[954]}), .bottom_right({trees[955], lumberyards[955]}), .init(2'b00), .state({trees[904], lumberyards[904]}));
acre acre_18_5 (.clk(clk), .en(en), .top_left({trees[854], lumberyards[854]}), .top({trees[855], lumberyards[855]}), .top_right({trees[856], lumberyards[856]}), .left({trees[904], lumberyards[904]}), .right({trees[906], lumberyards[906]}), .bottom_left({trees[954], lumberyards[954]}), .bottom({trees[955], lumberyards[955]}), .bottom_right({trees[956], lumberyards[956]}), .init(2'b00), .state({trees[905], lumberyards[905]}));
acre acre_18_6 (.clk(clk), .en(en), .top_left({trees[855], lumberyards[855]}), .top({trees[856], lumberyards[856]}), .top_right({trees[857], lumberyards[857]}), .left({trees[905], lumberyards[905]}), .right({trees[907], lumberyards[907]}), .bottom_left({trees[955], lumberyards[955]}), .bottom({trees[956], lumberyards[956]}), .bottom_right({trees[957], lumberyards[957]}), .init(2'b00), .state({trees[906], lumberyards[906]}));
acre acre_18_7 (.clk(clk), .en(en), .top_left({trees[856], lumberyards[856]}), .top({trees[857], lumberyards[857]}), .top_right({trees[858], lumberyards[858]}), .left({trees[906], lumberyards[906]}), .right({trees[908], lumberyards[908]}), .bottom_left({trees[956], lumberyards[956]}), .bottom({trees[957], lumberyards[957]}), .bottom_right({trees[958], lumberyards[958]}), .init(2'b00), .state({trees[907], lumberyards[907]}));
acre acre_18_8 (.clk(clk), .en(en), .top_left({trees[857], lumberyards[857]}), .top({trees[858], lumberyards[858]}), .top_right({trees[859], lumberyards[859]}), .left({trees[907], lumberyards[907]}), .right({trees[909], lumberyards[909]}), .bottom_left({trees[957], lumberyards[957]}), .bottom({trees[958], lumberyards[958]}), .bottom_right({trees[959], lumberyards[959]}), .init(2'b10), .state({trees[908], lumberyards[908]}));
acre acre_18_9 (.clk(clk), .en(en), .top_left({trees[858], lumberyards[858]}), .top({trees[859], lumberyards[859]}), .top_right({trees[860], lumberyards[860]}), .left({trees[908], lumberyards[908]}), .right({trees[910], lumberyards[910]}), .bottom_left({trees[958], lumberyards[958]}), .bottom({trees[959], lumberyards[959]}), .bottom_right({trees[960], lumberyards[960]}), .init(2'b00), .state({trees[909], lumberyards[909]}));
acre acre_18_10 (.clk(clk), .en(en), .top_left({trees[859], lumberyards[859]}), .top({trees[860], lumberyards[860]}), .top_right({trees[861], lumberyards[861]}), .left({trees[909], lumberyards[909]}), .right({trees[911], lumberyards[911]}), .bottom_left({trees[959], lumberyards[959]}), .bottom({trees[960], lumberyards[960]}), .bottom_right({trees[961], lumberyards[961]}), .init(2'b01), .state({trees[910], lumberyards[910]}));
acre acre_18_11 (.clk(clk), .en(en), .top_left({trees[860], lumberyards[860]}), .top({trees[861], lumberyards[861]}), .top_right({trees[862], lumberyards[862]}), .left({trees[910], lumberyards[910]}), .right({trees[912], lumberyards[912]}), .bottom_left({trees[960], lumberyards[960]}), .bottom({trees[961], lumberyards[961]}), .bottom_right({trees[962], lumberyards[962]}), .init(2'b01), .state({trees[911], lumberyards[911]}));
acre acre_18_12 (.clk(clk), .en(en), .top_left({trees[861], lumberyards[861]}), .top({trees[862], lumberyards[862]}), .top_right({trees[863], lumberyards[863]}), .left({trees[911], lumberyards[911]}), .right({trees[913], lumberyards[913]}), .bottom_left({trees[961], lumberyards[961]}), .bottom({trees[962], lumberyards[962]}), .bottom_right({trees[963], lumberyards[963]}), .init(2'b10), .state({trees[912], lumberyards[912]}));
acre acre_18_13 (.clk(clk), .en(en), .top_left({trees[862], lumberyards[862]}), .top({trees[863], lumberyards[863]}), .top_right({trees[864], lumberyards[864]}), .left({trees[912], lumberyards[912]}), .right({trees[914], lumberyards[914]}), .bottom_left({trees[962], lumberyards[962]}), .bottom({trees[963], lumberyards[963]}), .bottom_right({trees[964], lumberyards[964]}), .init(2'b00), .state({trees[913], lumberyards[913]}));
acre acre_18_14 (.clk(clk), .en(en), .top_left({trees[863], lumberyards[863]}), .top({trees[864], lumberyards[864]}), .top_right({trees[865], lumberyards[865]}), .left({trees[913], lumberyards[913]}), .right({trees[915], lumberyards[915]}), .bottom_left({trees[963], lumberyards[963]}), .bottom({trees[964], lumberyards[964]}), .bottom_right({trees[965], lumberyards[965]}), .init(2'b10), .state({trees[914], lumberyards[914]}));
acre acre_18_15 (.clk(clk), .en(en), .top_left({trees[864], lumberyards[864]}), .top({trees[865], lumberyards[865]}), .top_right({trees[866], lumberyards[866]}), .left({trees[914], lumberyards[914]}), .right({trees[916], lumberyards[916]}), .bottom_left({trees[964], lumberyards[964]}), .bottom({trees[965], lumberyards[965]}), .bottom_right({trees[966], lumberyards[966]}), .init(2'b10), .state({trees[915], lumberyards[915]}));
acre acre_18_16 (.clk(clk), .en(en), .top_left({trees[865], lumberyards[865]}), .top({trees[866], lumberyards[866]}), .top_right({trees[867], lumberyards[867]}), .left({trees[915], lumberyards[915]}), .right({trees[917], lumberyards[917]}), .bottom_left({trees[965], lumberyards[965]}), .bottom({trees[966], lumberyards[966]}), .bottom_right({trees[967], lumberyards[967]}), .init(2'b00), .state({trees[916], lumberyards[916]}));
acre acre_18_17 (.clk(clk), .en(en), .top_left({trees[866], lumberyards[866]}), .top({trees[867], lumberyards[867]}), .top_right({trees[868], lumberyards[868]}), .left({trees[916], lumberyards[916]}), .right({trees[918], lumberyards[918]}), .bottom_left({trees[966], lumberyards[966]}), .bottom({trees[967], lumberyards[967]}), .bottom_right({trees[968], lumberyards[968]}), .init(2'b00), .state({trees[917], lumberyards[917]}));
acre acre_18_18 (.clk(clk), .en(en), .top_left({trees[867], lumberyards[867]}), .top({trees[868], lumberyards[868]}), .top_right({trees[869], lumberyards[869]}), .left({trees[917], lumberyards[917]}), .right({trees[919], lumberyards[919]}), .bottom_left({trees[967], lumberyards[967]}), .bottom({trees[968], lumberyards[968]}), .bottom_right({trees[969], lumberyards[969]}), .init(2'b01), .state({trees[918], lumberyards[918]}));
acre acre_18_19 (.clk(clk), .en(en), .top_left({trees[868], lumberyards[868]}), .top({trees[869], lumberyards[869]}), .top_right({trees[870], lumberyards[870]}), .left({trees[918], lumberyards[918]}), .right({trees[920], lumberyards[920]}), .bottom_left({trees[968], lumberyards[968]}), .bottom({trees[969], lumberyards[969]}), .bottom_right({trees[970], lumberyards[970]}), .init(2'b10), .state({trees[919], lumberyards[919]}));
acre acre_18_20 (.clk(clk), .en(en), .top_left({trees[869], lumberyards[869]}), .top({trees[870], lumberyards[870]}), .top_right({trees[871], lumberyards[871]}), .left({trees[919], lumberyards[919]}), .right({trees[921], lumberyards[921]}), .bottom_left({trees[969], lumberyards[969]}), .bottom({trees[970], lumberyards[970]}), .bottom_right({trees[971], lumberyards[971]}), .init(2'b10), .state({trees[920], lumberyards[920]}));
acre acre_18_21 (.clk(clk), .en(en), .top_left({trees[870], lumberyards[870]}), .top({trees[871], lumberyards[871]}), .top_right({trees[872], lumberyards[872]}), .left({trees[920], lumberyards[920]}), .right({trees[922], lumberyards[922]}), .bottom_left({trees[970], lumberyards[970]}), .bottom({trees[971], lumberyards[971]}), .bottom_right({trees[972], lumberyards[972]}), .init(2'b00), .state({trees[921], lumberyards[921]}));
acre acre_18_22 (.clk(clk), .en(en), .top_left({trees[871], lumberyards[871]}), .top({trees[872], lumberyards[872]}), .top_right({trees[873], lumberyards[873]}), .left({trees[921], lumberyards[921]}), .right({trees[923], lumberyards[923]}), .bottom_left({trees[971], lumberyards[971]}), .bottom({trees[972], lumberyards[972]}), .bottom_right({trees[973], lumberyards[973]}), .init(2'b10), .state({trees[922], lumberyards[922]}));
acre acre_18_23 (.clk(clk), .en(en), .top_left({trees[872], lumberyards[872]}), .top({trees[873], lumberyards[873]}), .top_right({trees[874], lumberyards[874]}), .left({trees[922], lumberyards[922]}), .right({trees[924], lumberyards[924]}), .bottom_left({trees[972], lumberyards[972]}), .bottom({trees[973], lumberyards[973]}), .bottom_right({trees[974], lumberyards[974]}), .init(2'b01), .state({trees[923], lumberyards[923]}));
acre acre_18_24 (.clk(clk), .en(en), .top_left({trees[873], lumberyards[873]}), .top({trees[874], lumberyards[874]}), .top_right({trees[875], lumberyards[875]}), .left({trees[923], lumberyards[923]}), .right({trees[925], lumberyards[925]}), .bottom_left({trees[973], lumberyards[973]}), .bottom({trees[974], lumberyards[974]}), .bottom_right({trees[975], lumberyards[975]}), .init(2'b10), .state({trees[924], lumberyards[924]}));
acre acre_18_25 (.clk(clk), .en(en), .top_left({trees[874], lumberyards[874]}), .top({trees[875], lumberyards[875]}), .top_right({trees[876], lumberyards[876]}), .left({trees[924], lumberyards[924]}), .right({trees[926], lumberyards[926]}), .bottom_left({trees[974], lumberyards[974]}), .bottom({trees[975], lumberyards[975]}), .bottom_right({trees[976], lumberyards[976]}), .init(2'b00), .state({trees[925], lumberyards[925]}));
acre acre_18_26 (.clk(clk), .en(en), .top_left({trees[875], lumberyards[875]}), .top({trees[876], lumberyards[876]}), .top_right({trees[877], lumberyards[877]}), .left({trees[925], lumberyards[925]}), .right({trees[927], lumberyards[927]}), .bottom_left({trees[975], lumberyards[975]}), .bottom({trees[976], lumberyards[976]}), .bottom_right({trees[977], lumberyards[977]}), .init(2'b00), .state({trees[926], lumberyards[926]}));
acre acre_18_27 (.clk(clk), .en(en), .top_left({trees[876], lumberyards[876]}), .top({trees[877], lumberyards[877]}), .top_right({trees[878], lumberyards[878]}), .left({trees[926], lumberyards[926]}), .right({trees[928], lumberyards[928]}), .bottom_left({trees[976], lumberyards[976]}), .bottom({trees[977], lumberyards[977]}), .bottom_right({trees[978], lumberyards[978]}), .init(2'b00), .state({trees[927], lumberyards[927]}));
acre acre_18_28 (.clk(clk), .en(en), .top_left({trees[877], lumberyards[877]}), .top({trees[878], lumberyards[878]}), .top_right({trees[879], lumberyards[879]}), .left({trees[927], lumberyards[927]}), .right({trees[929], lumberyards[929]}), .bottom_left({trees[977], lumberyards[977]}), .bottom({trees[978], lumberyards[978]}), .bottom_right({trees[979], lumberyards[979]}), .init(2'b01), .state({trees[928], lumberyards[928]}));
acre acre_18_29 (.clk(clk), .en(en), .top_left({trees[878], lumberyards[878]}), .top({trees[879], lumberyards[879]}), .top_right({trees[880], lumberyards[880]}), .left({trees[928], lumberyards[928]}), .right({trees[930], lumberyards[930]}), .bottom_left({trees[978], lumberyards[978]}), .bottom({trees[979], lumberyards[979]}), .bottom_right({trees[980], lumberyards[980]}), .init(2'b00), .state({trees[929], lumberyards[929]}));
acre acre_18_30 (.clk(clk), .en(en), .top_left({trees[879], lumberyards[879]}), .top({trees[880], lumberyards[880]}), .top_right({trees[881], lumberyards[881]}), .left({trees[929], lumberyards[929]}), .right({trees[931], lumberyards[931]}), .bottom_left({trees[979], lumberyards[979]}), .bottom({trees[980], lumberyards[980]}), .bottom_right({trees[981], lumberyards[981]}), .init(2'b00), .state({trees[930], lumberyards[930]}));
acre acre_18_31 (.clk(clk), .en(en), .top_left({trees[880], lumberyards[880]}), .top({trees[881], lumberyards[881]}), .top_right({trees[882], lumberyards[882]}), .left({trees[930], lumberyards[930]}), .right({trees[932], lumberyards[932]}), .bottom_left({trees[980], lumberyards[980]}), .bottom({trees[981], lumberyards[981]}), .bottom_right({trees[982], lumberyards[982]}), .init(2'b01), .state({trees[931], lumberyards[931]}));
acre acre_18_32 (.clk(clk), .en(en), .top_left({trees[881], lumberyards[881]}), .top({trees[882], lumberyards[882]}), .top_right({trees[883], lumberyards[883]}), .left({trees[931], lumberyards[931]}), .right({trees[933], lumberyards[933]}), .bottom_left({trees[981], lumberyards[981]}), .bottom({trees[982], lumberyards[982]}), .bottom_right({trees[983], lumberyards[983]}), .init(2'b10), .state({trees[932], lumberyards[932]}));
acre acre_18_33 (.clk(clk), .en(en), .top_left({trees[882], lumberyards[882]}), .top({trees[883], lumberyards[883]}), .top_right({trees[884], lumberyards[884]}), .left({trees[932], lumberyards[932]}), .right({trees[934], lumberyards[934]}), .bottom_left({trees[982], lumberyards[982]}), .bottom({trees[983], lumberyards[983]}), .bottom_right({trees[984], lumberyards[984]}), .init(2'b01), .state({trees[933], lumberyards[933]}));
acre acre_18_34 (.clk(clk), .en(en), .top_left({trees[883], lumberyards[883]}), .top({trees[884], lumberyards[884]}), .top_right({trees[885], lumberyards[885]}), .left({trees[933], lumberyards[933]}), .right({trees[935], lumberyards[935]}), .bottom_left({trees[983], lumberyards[983]}), .bottom({trees[984], lumberyards[984]}), .bottom_right({trees[985], lumberyards[985]}), .init(2'b10), .state({trees[934], lumberyards[934]}));
acre acre_18_35 (.clk(clk), .en(en), .top_left({trees[884], lumberyards[884]}), .top({trees[885], lumberyards[885]}), .top_right({trees[886], lumberyards[886]}), .left({trees[934], lumberyards[934]}), .right({trees[936], lumberyards[936]}), .bottom_left({trees[984], lumberyards[984]}), .bottom({trees[985], lumberyards[985]}), .bottom_right({trees[986], lumberyards[986]}), .init(2'b00), .state({trees[935], lumberyards[935]}));
acre acre_18_36 (.clk(clk), .en(en), .top_left({trees[885], lumberyards[885]}), .top({trees[886], lumberyards[886]}), .top_right({trees[887], lumberyards[887]}), .left({trees[935], lumberyards[935]}), .right({trees[937], lumberyards[937]}), .bottom_left({trees[985], lumberyards[985]}), .bottom({trees[986], lumberyards[986]}), .bottom_right({trees[987], lumberyards[987]}), .init(2'b01), .state({trees[936], lumberyards[936]}));
acre acre_18_37 (.clk(clk), .en(en), .top_left({trees[886], lumberyards[886]}), .top({trees[887], lumberyards[887]}), .top_right({trees[888], lumberyards[888]}), .left({trees[936], lumberyards[936]}), .right({trees[938], lumberyards[938]}), .bottom_left({trees[986], lumberyards[986]}), .bottom({trees[987], lumberyards[987]}), .bottom_right({trees[988], lumberyards[988]}), .init(2'b00), .state({trees[937], lumberyards[937]}));
acre acre_18_38 (.clk(clk), .en(en), .top_left({trees[887], lumberyards[887]}), .top({trees[888], lumberyards[888]}), .top_right({trees[889], lumberyards[889]}), .left({trees[937], lumberyards[937]}), .right({trees[939], lumberyards[939]}), .bottom_left({trees[987], lumberyards[987]}), .bottom({trees[988], lumberyards[988]}), .bottom_right({trees[989], lumberyards[989]}), .init(2'b10), .state({trees[938], lumberyards[938]}));
acre acre_18_39 (.clk(clk), .en(en), .top_left({trees[888], lumberyards[888]}), .top({trees[889], lumberyards[889]}), .top_right({trees[890], lumberyards[890]}), .left({trees[938], lumberyards[938]}), .right({trees[940], lumberyards[940]}), .bottom_left({trees[988], lumberyards[988]}), .bottom({trees[989], lumberyards[989]}), .bottom_right({trees[990], lumberyards[990]}), .init(2'b00), .state({trees[939], lumberyards[939]}));
acre acre_18_40 (.clk(clk), .en(en), .top_left({trees[889], lumberyards[889]}), .top({trees[890], lumberyards[890]}), .top_right({trees[891], lumberyards[891]}), .left({trees[939], lumberyards[939]}), .right({trees[941], lumberyards[941]}), .bottom_left({trees[989], lumberyards[989]}), .bottom({trees[990], lumberyards[990]}), .bottom_right({trees[991], lumberyards[991]}), .init(2'b01), .state({trees[940], lumberyards[940]}));
acre acre_18_41 (.clk(clk), .en(en), .top_left({trees[890], lumberyards[890]}), .top({trees[891], lumberyards[891]}), .top_right({trees[892], lumberyards[892]}), .left({trees[940], lumberyards[940]}), .right({trees[942], lumberyards[942]}), .bottom_left({trees[990], lumberyards[990]}), .bottom({trees[991], lumberyards[991]}), .bottom_right({trees[992], lumberyards[992]}), .init(2'b00), .state({trees[941], lumberyards[941]}));
acre acre_18_42 (.clk(clk), .en(en), .top_left({trees[891], lumberyards[891]}), .top({trees[892], lumberyards[892]}), .top_right({trees[893], lumberyards[893]}), .left({trees[941], lumberyards[941]}), .right({trees[943], lumberyards[943]}), .bottom_left({trees[991], lumberyards[991]}), .bottom({trees[992], lumberyards[992]}), .bottom_right({trees[993], lumberyards[993]}), .init(2'b00), .state({trees[942], lumberyards[942]}));
acre acre_18_43 (.clk(clk), .en(en), .top_left({trees[892], lumberyards[892]}), .top({trees[893], lumberyards[893]}), .top_right({trees[894], lumberyards[894]}), .left({trees[942], lumberyards[942]}), .right({trees[944], lumberyards[944]}), .bottom_left({trees[992], lumberyards[992]}), .bottom({trees[993], lumberyards[993]}), .bottom_right({trees[994], lumberyards[994]}), .init(2'b00), .state({trees[943], lumberyards[943]}));
acre acre_18_44 (.clk(clk), .en(en), .top_left({trees[893], lumberyards[893]}), .top({trees[894], lumberyards[894]}), .top_right({trees[895], lumberyards[895]}), .left({trees[943], lumberyards[943]}), .right({trees[945], lumberyards[945]}), .bottom_left({trees[993], lumberyards[993]}), .bottom({trees[994], lumberyards[994]}), .bottom_right({trees[995], lumberyards[995]}), .init(2'b00), .state({trees[944], lumberyards[944]}));
acre acre_18_45 (.clk(clk), .en(en), .top_left({trees[894], lumberyards[894]}), .top({trees[895], lumberyards[895]}), .top_right({trees[896], lumberyards[896]}), .left({trees[944], lumberyards[944]}), .right({trees[946], lumberyards[946]}), .bottom_left({trees[994], lumberyards[994]}), .bottom({trees[995], lumberyards[995]}), .bottom_right({trees[996], lumberyards[996]}), .init(2'b00), .state({trees[945], lumberyards[945]}));
acre acre_18_46 (.clk(clk), .en(en), .top_left({trees[895], lumberyards[895]}), .top({trees[896], lumberyards[896]}), .top_right({trees[897], lumberyards[897]}), .left({trees[945], lumberyards[945]}), .right({trees[947], lumberyards[947]}), .bottom_left({trees[995], lumberyards[995]}), .bottom({trees[996], lumberyards[996]}), .bottom_right({trees[997], lumberyards[997]}), .init(2'b00), .state({trees[946], lumberyards[946]}));
acre acre_18_47 (.clk(clk), .en(en), .top_left({trees[896], lumberyards[896]}), .top({trees[897], lumberyards[897]}), .top_right({trees[898], lumberyards[898]}), .left({trees[946], lumberyards[946]}), .right({trees[948], lumberyards[948]}), .bottom_left({trees[996], lumberyards[996]}), .bottom({trees[997], lumberyards[997]}), .bottom_right({trees[998], lumberyards[998]}), .init(2'b00), .state({trees[947], lumberyards[947]}));
acre acre_18_48 (.clk(clk), .en(en), .top_left({trees[897], lumberyards[897]}), .top({trees[898], lumberyards[898]}), .top_right({trees[899], lumberyards[899]}), .left({trees[947], lumberyards[947]}), .right({trees[949], lumberyards[949]}), .bottom_left({trees[997], lumberyards[997]}), .bottom({trees[998], lumberyards[998]}), .bottom_right({trees[999], lumberyards[999]}), .init(2'b00), .state({trees[948], lumberyards[948]}));
acre acre_18_49 (.clk(clk), .en(en), .top_left({trees[898], lumberyards[898]}), .top({trees[899], lumberyards[899]}), .top_right(2'b0), .left({trees[948], lumberyards[948]}), .right(2'b0), .bottom_left({trees[998], lumberyards[998]}), .bottom({trees[999], lumberyards[999]}), .bottom_right(2'b0), .init(2'b01), .state({trees[949], lumberyards[949]}));
acre acre_19_0 (.clk(clk), .en(en), .top_left(2'b0), .top({trees[900], lumberyards[900]}), .top_right({trees[901], lumberyards[901]}), .left(2'b0), .right({trees[951], lumberyards[951]}), .bottom_left(2'b0), .bottom({trees[1000], lumberyards[1000]}), .bottom_right({trees[1001], lumberyards[1001]}), .init(2'b01), .state({trees[950], lumberyards[950]}));
acre acre_19_1 (.clk(clk), .en(en), .top_left({trees[900], lumberyards[900]}), .top({trees[901], lumberyards[901]}), .top_right({trees[902], lumberyards[902]}), .left({trees[950], lumberyards[950]}), .right({trees[952], lumberyards[952]}), .bottom_left({trees[1000], lumberyards[1000]}), .bottom({trees[1001], lumberyards[1001]}), .bottom_right({trees[1002], lumberyards[1002]}), .init(2'b00), .state({trees[951], lumberyards[951]}));
acre acre_19_2 (.clk(clk), .en(en), .top_left({trees[901], lumberyards[901]}), .top({trees[902], lumberyards[902]}), .top_right({trees[903], lumberyards[903]}), .left({trees[951], lumberyards[951]}), .right({trees[953], lumberyards[953]}), .bottom_left({trees[1001], lumberyards[1001]}), .bottom({trees[1002], lumberyards[1002]}), .bottom_right({trees[1003], lumberyards[1003]}), .init(2'b10), .state({trees[952], lumberyards[952]}));
acre acre_19_3 (.clk(clk), .en(en), .top_left({trees[902], lumberyards[902]}), .top({trees[903], lumberyards[903]}), .top_right({trees[904], lumberyards[904]}), .left({trees[952], lumberyards[952]}), .right({trees[954], lumberyards[954]}), .bottom_left({trees[1002], lumberyards[1002]}), .bottom({trees[1003], lumberyards[1003]}), .bottom_right({trees[1004], lumberyards[1004]}), .init(2'b00), .state({trees[953], lumberyards[953]}));
acre acre_19_4 (.clk(clk), .en(en), .top_left({trees[903], lumberyards[903]}), .top({trees[904], lumberyards[904]}), .top_right({trees[905], lumberyards[905]}), .left({trees[953], lumberyards[953]}), .right({trees[955], lumberyards[955]}), .bottom_left({trees[1003], lumberyards[1003]}), .bottom({trees[1004], lumberyards[1004]}), .bottom_right({trees[1005], lumberyards[1005]}), .init(2'b10), .state({trees[954], lumberyards[954]}));
acre acre_19_5 (.clk(clk), .en(en), .top_left({trees[904], lumberyards[904]}), .top({trees[905], lumberyards[905]}), .top_right({trees[906], lumberyards[906]}), .left({trees[954], lumberyards[954]}), .right({trees[956], lumberyards[956]}), .bottom_left({trees[1004], lumberyards[1004]}), .bottom({trees[1005], lumberyards[1005]}), .bottom_right({trees[1006], lumberyards[1006]}), .init(2'b10), .state({trees[955], lumberyards[955]}));
acre acre_19_6 (.clk(clk), .en(en), .top_left({trees[905], lumberyards[905]}), .top({trees[906], lumberyards[906]}), .top_right({trees[907], lumberyards[907]}), .left({trees[955], lumberyards[955]}), .right({trees[957], lumberyards[957]}), .bottom_left({trees[1005], lumberyards[1005]}), .bottom({trees[1006], lumberyards[1006]}), .bottom_right({trees[1007], lumberyards[1007]}), .init(2'b00), .state({trees[956], lumberyards[956]}));
acre acre_19_7 (.clk(clk), .en(en), .top_left({trees[906], lumberyards[906]}), .top({trees[907], lumberyards[907]}), .top_right({trees[908], lumberyards[908]}), .left({trees[956], lumberyards[956]}), .right({trees[958], lumberyards[958]}), .bottom_left({trees[1006], lumberyards[1006]}), .bottom({trees[1007], lumberyards[1007]}), .bottom_right({trees[1008], lumberyards[1008]}), .init(2'b00), .state({trees[957], lumberyards[957]}));
acre acre_19_8 (.clk(clk), .en(en), .top_left({trees[907], lumberyards[907]}), .top({trees[908], lumberyards[908]}), .top_right({trees[909], lumberyards[909]}), .left({trees[957], lumberyards[957]}), .right({trees[959], lumberyards[959]}), .bottom_left({trees[1007], lumberyards[1007]}), .bottom({trees[1008], lumberyards[1008]}), .bottom_right({trees[1009], lumberyards[1009]}), .init(2'b10), .state({trees[958], lumberyards[958]}));
acre acre_19_9 (.clk(clk), .en(en), .top_left({trees[908], lumberyards[908]}), .top({trees[909], lumberyards[909]}), .top_right({trees[910], lumberyards[910]}), .left({trees[958], lumberyards[958]}), .right({trees[960], lumberyards[960]}), .bottom_left({trees[1008], lumberyards[1008]}), .bottom({trees[1009], lumberyards[1009]}), .bottom_right({trees[1010], lumberyards[1010]}), .init(2'b10), .state({trees[959], lumberyards[959]}));
acre acre_19_10 (.clk(clk), .en(en), .top_left({trees[909], lumberyards[909]}), .top({trees[910], lumberyards[910]}), .top_right({trees[911], lumberyards[911]}), .left({trees[959], lumberyards[959]}), .right({trees[961], lumberyards[961]}), .bottom_left({trees[1009], lumberyards[1009]}), .bottom({trees[1010], lumberyards[1010]}), .bottom_right({trees[1011], lumberyards[1011]}), .init(2'b00), .state({trees[960], lumberyards[960]}));
acre acre_19_11 (.clk(clk), .en(en), .top_left({trees[910], lumberyards[910]}), .top({trees[911], lumberyards[911]}), .top_right({trees[912], lumberyards[912]}), .left({trees[960], lumberyards[960]}), .right({trees[962], lumberyards[962]}), .bottom_left({trees[1010], lumberyards[1010]}), .bottom({trees[1011], lumberyards[1011]}), .bottom_right({trees[1012], lumberyards[1012]}), .init(2'b01), .state({trees[961], lumberyards[961]}));
acre acre_19_12 (.clk(clk), .en(en), .top_left({trees[911], lumberyards[911]}), .top({trees[912], lumberyards[912]}), .top_right({trees[913], lumberyards[913]}), .left({trees[961], lumberyards[961]}), .right({trees[963], lumberyards[963]}), .bottom_left({trees[1011], lumberyards[1011]}), .bottom({trees[1012], lumberyards[1012]}), .bottom_right({trees[1013], lumberyards[1013]}), .init(2'b00), .state({trees[962], lumberyards[962]}));
acre acre_19_13 (.clk(clk), .en(en), .top_left({trees[912], lumberyards[912]}), .top({trees[913], lumberyards[913]}), .top_right({trees[914], lumberyards[914]}), .left({trees[962], lumberyards[962]}), .right({trees[964], lumberyards[964]}), .bottom_left({trees[1012], lumberyards[1012]}), .bottom({trees[1013], lumberyards[1013]}), .bottom_right({trees[1014], lumberyards[1014]}), .init(2'b00), .state({trees[963], lumberyards[963]}));
acre acre_19_14 (.clk(clk), .en(en), .top_left({trees[913], lumberyards[913]}), .top({trees[914], lumberyards[914]}), .top_right({trees[915], lumberyards[915]}), .left({trees[963], lumberyards[963]}), .right({trees[965], lumberyards[965]}), .bottom_left({trees[1013], lumberyards[1013]}), .bottom({trees[1014], lumberyards[1014]}), .bottom_right({trees[1015], lumberyards[1015]}), .init(2'b00), .state({trees[964], lumberyards[964]}));
acre acre_19_15 (.clk(clk), .en(en), .top_left({trees[914], lumberyards[914]}), .top({trees[915], lumberyards[915]}), .top_right({trees[916], lumberyards[916]}), .left({trees[964], lumberyards[964]}), .right({trees[966], lumberyards[966]}), .bottom_left({trees[1014], lumberyards[1014]}), .bottom({trees[1015], lumberyards[1015]}), .bottom_right({trees[1016], lumberyards[1016]}), .init(2'b10), .state({trees[965], lumberyards[965]}));
acre acre_19_16 (.clk(clk), .en(en), .top_left({trees[915], lumberyards[915]}), .top({trees[916], lumberyards[916]}), .top_right({trees[917], lumberyards[917]}), .left({trees[965], lumberyards[965]}), .right({trees[967], lumberyards[967]}), .bottom_left({trees[1015], lumberyards[1015]}), .bottom({trees[1016], lumberyards[1016]}), .bottom_right({trees[1017], lumberyards[1017]}), .init(2'b10), .state({trees[966], lumberyards[966]}));
acre acre_19_17 (.clk(clk), .en(en), .top_left({trees[916], lumberyards[916]}), .top({trees[917], lumberyards[917]}), .top_right({trees[918], lumberyards[918]}), .left({trees[966], lumberyards[966]}), .right({trees[968], lumberyards[968]}), .bottom_left({trees[1016], lumberyards[1016]}), .bottom({trees[1017], lumberyards[1017]}), .bottom_right({trees[1018], lumberyards[1018]}), .init(2'b00), .state({trees[967], lumberyards[967]}));
acre acre_19_18 (.clk(clk), .en(en), .top_left({trees[917], lumberyards[917]}), .top({trees[918], lumberyards[918]}), .top_right({trees[919], lumberyards[919]}), .left({trees[967], lumberyards[967]}), .right({trees[969], lumberyards[969]}), .bottom_left({trees[1017], lumberyards[1017]}), .bottom({trees[1018], lumberyards[1018]}), .bottom_right({trees[1019], lumberyards[1019]}), .init(2'b00), .state({trees[968], lumberyards[968]}));
acre acre_19_19 (.clk(clk), .en(en), .top_left({trees[918], lumberyards[918]}), .top({trees[919], lumberyards[919]}), .top_right({trees[920], lumberyards[920]}), .left({trees[968], lumberyards[968]}), .right({trees[970], lumberyards[970]}), .bottom_left({trees[1018], lumberyards[1018]}), .bottom({trees[1019], lumberyards[1019]}), .bottom_right({trees[1020], lumberyards[1020]}), .init(2'b01), .state({trees[969], lumberyards[969]}));
acre acre_19_20 (.clk(clk), .en(en), .top_left({trees[919], lumberyards[919]}), .top({trees[920], lumberyards[920]}), .top_right({trees[921], lumberyards[921]}), .left({trees[969], lumberyards[969]}), .right({trees[971], lumberyards[971]}), .bottom_left({trees[1019], lumberyards[1019]}), .bottom({trees[1020], lumberyards[1020]}), .bottom_right({trees[1021], lumberyards[1021]}), .init(2'b01), .state({trees[970], lumberyards[970]}));
acre acre_19_21 (.clk(clk), .en(en), .top_left({trees[920], lumberyards[920]}), .top({trees[921], lumberyards[921]}), .top_right({trees[922], lumberyards[922]}), .left({trees[970], lumberyards[970]}), .right({trees[972], lumberyards[972]}), .bottom_left({trees[1020], lumberyards[1020]}), .bottom({trees[1021], lumberyards[1021]}), .bottom_right({trees[1022], lumberyards[1022]}), .init(2'b00), .state({trees[971], lumberyards[971]}));
acre acre_19_22 (.clk(clk), .en(en), .top_left({trees[921], lumberyards[921]}), .top({trees[922], lumberyards[922]}), .top_right({trees[923], lumberyards[923]}), .left({trees[971], lumberyards[971]}), .right({trees[973], lumberyards[973]}), .bottom_left({trees[1021], lumberyards[1021]}), .bottom({trees[1022], lumberyards[1022]}), .bottom_right({trees[1023], lumberyards[1023]}), .init(2'b00), .state({trees[972], lumberyards[972]}));
acre acre_19_23 (.clk(clk), .en(en), .top_left({trees[922], lumberyards[922]}), .top({trees[923], lumberyards[923]}), .top_right({trees[924], lumberyards[924]}), .left({trees[972], lumberyards[972]}), .right({trees[974], lumberyards[974]}), .bottom_left({trees[1022], lumberyards[1022]}), .bottom({trees[1023], lumberyards[1023]}), .bottom_right({trees[1024], lumberyards[1024]}), .init(2'b10), .state({trees[973], lumberyards[973]}));
acre acre_19_24 (.clk(clk), .en(en), .top_left({trees[923], lumberyards[923]}), .top({trees[924], lumberyards[924]}), .top_right({trees[925], lumberyards[925]}), .left({trees[973], lumberyards[973]}), .right({trees[975], lumberyards[975]}), .bottom_left({trees[1023], lumberyards[1023]}), .bottom({trees[1024], lumberyards[1024]}), .bottom_right({trees[1025], lumberyards[1025]}), .init(2'b01), .state({trees[974], lumberyards[974]}));
acre acre_19_25 (.clk(clk), .en(en), .top_left({trees[924], lumberyards[924]}), .top({trees[925], lumberyards[925]}), .top_right({trees[926], lumberyards[926]}), .left({trees[974], lumberyards[974]}), .right({trees[976], lumberyards[976]}), .bottom_left({trees[1024], lumberyards[1024]}), .bottom({trees[1025], lumberyards[1025]}), .bottom_right({trees[1026], lumberyards[1026]}), .init(2'b00), .state({trees[975], lumberyards[975]}));
acre acre_19_26 (.clk(clk), .en(en), .top_left({trees[925], lumberyards[925]}), .top({trees[926], lumberyards[926]}), .top_right({trees[927], lumberyards[927]}), .left({trees[975], lumberyards[975]}), .right({trees[977], lumberyards[977]}), .bottom_left({trees[1025], lumberyards[1025]}), .bottom({trees[1026], lumberyards[1026]}), .bottom_right({trees[1027], lumberyards[1027]}), .init(2'b00), .state({trees[976], lumberyards[976]}));
acre acre_19_27 (.clk(clk), .en(en), .top_left({trees[926], lumberyards[926]}), .top({trees[927], lumberyards[927]}), .top_right({trees[928], lumberyards[928]}), .left({trees[976], lumberyards[976]}), .right({trees[978], lumberyards[978]}), .bottom_left({trees[1026], lumberyards[1026]}), .bottom({trees[1027], lumberyards[1027]}), .bottom_right({trees[1028], lumberyards[1028]}), .init(2'b00), .state({trees[977], lumberyards[977]}));
acre acre_19_28 (.clk(clk), .en(en), .top_left({trees[927], lumberyards[927]}), .top({trees[928], lumberyards[928]}), .top_right({trees[929], lumberyards[929]}), .left({trees[977], lumberyards[977]}), .right({trees[979], lumberyards[979]}), .bottom_left({trees[1027], lumberyards[1027]}), .bottom({trees[1028], lumberyards[1028]}), .bottom_right({trees[1029], lumberyards[1029]}), .init(2'b00), .state({trees[978], lumberyards[978]}));
acre acre_19_29 (.clk(clk), .en(en), .top_left({trees[928], lumberyards[928]}), .top({trees[929], lumberyards[929]}), .top_right({trees[930], lumberyards[930]}), .left({trees[978], lumberyards[978]}), .right({trees[980], lumberyards[980]}), .bottom_left({trees[1028], lumberyards[1028]}), .bottom({trees[1029], lumberyards[1029]}), .bottom_right({trees[1030], lumberyards[1030]}), .init(2'b01), .state({trees[979], lumberyards[979]}));
acre acre_19_30 (.clk(clk), .en(en), .top_left({trees[929], lumberyards[929]}), .top({trees[930], lumberyards[930]}), .top_right({trees[931], lumberyards[931]}), .left({trees[979], lumberyards[979]}), .right({trees[981], lumberyards[981]}), .bottom_left({trees[1029], lumberyards[1029]}), .bottom({trees[1030], lumberyards[1030]}), .bottom_right({trees[1031], lumberyards[1031]}), .init(2'b10), .state({trees[980], lumberyards[980]}));
acre acre_19_31 (.clk(clk), .en(en), .top_left({trees[930], lumberyards[930]}), .top({trees[931], lumberyards[931]}), .top_right({trees[932], lumberyards[932]}), .left({trees[980], lumberyards[980]}), .right({trees[982], lumberyards[982]}), .bottom_left({trees[1030], lumberyards[1030]}), .bottom({trees[1031], lumberyards[1031]}), .bottom_right({trees[1032], lumberyards[1032]}), .init(2'b00), .state({trees[981], lumberyards[981]}));
acre acre_19_32 (.clk(clk), .en(en), .top_left({trees[931], lumberyards[931]}), .top({trees[932], lumberyards[932]}), .top_right({trees[933], lumberyards[933]}), .left({trees[981], lumberyards[981]}), .right({trees[983], lumberyards[983]}), .bottom_left({trees[1031], lumberyards[1031]}), .bottom({trees[1032], lumberyards[1032]}), .bottom_right({trees[1033], lumberyards[1033]}), .init(2'b00), .state({trees[982], lumberyards[982]}));
acre acre_19_33 (.clk(clk), .en(en), .top_left({trees[932], lumberyards[932]}), .top({trees[933], lumberyards[933]}), .top_right({trees[934], lumberyards[934]}), .left({trees[982], lumberyards[982]}), .right({trees[984], lumberyards[984]}), .bottom_left({trees[1032], lumberyards[1032]}), .bottom({trees[1033], lumberyards[1033]}), .bottom_right({trees[1034], lumberyards[1034]}), .init(2'b00), .state({trees[983], lumberyards[983]}));
acre acre_19_34 (.clk(clk), .en(en), .top_left({trees[933], lumberyards[933]}), .top({trees[934], lumberyards[934]}), .top_right({trees[935], lumberyards[935]}), .left({trees[983], lumberyards[983]}), .right({trees[985], lumberyards[985]}), .bottom_left({trees[1033], lumberyards[1033]}), .bottom({trees[1034], lumberyards[1034]}), .bottom_right({trees[1035], lumberyards[1035]}), .init(2'b00), .state({trees[984], lumberyards[984]}));
acre acre_19_35 (.clk(clk), .en(en), .top_left({trees[934], lumberyards[934]}), .top({trees[935], lumberyards[935]}), .top_right({trees[936], lumberyards[936]}), .left({trees[984], lumberyards[984]}), .right({trees[986], lumberyards[986]}), .bottom_left({trees[1034], lumberyards[1034]}), .bottom({trees[1035], lumberyards[1035]}), .bottom_right({trees[1036], lumberyards[1036]}), .init(2'b00), .state({trees[985], lumberyards[985]}));
acre acre_19_36 (.clk(clk), .en(en), .top_left({trees[935], lumberyards[935]}), .top({trees[936], lumberyards[936]}), .top_right({trees[937], lumberyards[937]}), .left({trees[985], lumberyards[985]}), .right({trees[987], lumberyards[987]}), .bottom_left({trees[1035], lumberyards[1035]}), .bottom({trees[1036], lumberyards[1036]}), .bottom_right({trees[1037], lumberyards[1037]}), .init(2'b10), .state({trees[986], lumberyards[986]}));
acre acre_19_37 (.clk(clk), .en(en), .top_left({trees[936], lumberyards[936]}), .top({trees[937], lumberyards[937]}), .top_right({trees[938], lumberyards[938]}), .left({trees[986], lumberyards[986]}), .right({trees[988], lumberyards[988]}), .bottom_left({trees[1036], lumberyards[1036]}), .bottom({trees[1037], lumberyards[1037]}), .bottom_right({trees[1038], lumberyards[1038]}), .init(2'b00), .state({trees[987], lumberyards[987]}));
acre acre_19_38 (.clk(clk), .en(en), .top_left({trees[937], lumberyards[937]}), .top({trees[938], lumberyards[938]}), .top_right({trees[939], lumberyards[939]}), .left({trees[987], lumberyards[987]}), .right({trees[989], lumberyards[989]}), .bottom_left({trees[1037], lumberyards[1037]}), .bottom({trees[1038], lumberyards[1038]}), .bottom_right({trees[1039], lumberyards[1039]}), .init(2'b00), .state({trees[988], lumberyards[988]}));
acre acre_19_39 (.clk(clk), .en(en), .top_left({trees[938], lumberyards[938]}), .top({trees[939], lumberyards[939]}), .top_right({trees[940], lumberyards[940]}), .left({trees[988], lumberyards[988]}), .right({trees[990], lumberyards[990]}), .bottom_left({trees[1038], lumberyards[1038]}), .bottom({trees[1039], lumberyards[1039]}), .bottom_right({trees[1040], lumberyards[1040]}), .init(2'b01), .state({trees[989], lumberyards[989]}));
acre acre_19_40 (.clk(clk), .en(en), .top_left({trees[939], lumberyards[939]}), .top({trees[940], lumberyards[940]}), .top_right({trees[941], lumberyards[941]}), .left({trees[989], lumberyards[989]}), .right({trees[991], lumberyards[991]}), .bottom_left({trees[1039], lumberyards[1039]}), .bottom({trees[1040], lumberyards[1040]}), .bottom_right({trees[1041], lumberyards[1041]}), .init(2'b00), .state({trees[990], lumberyards[990]}));
acre acre_19_41 (.clk(clk), .en(en), .top_left({trees[940], lumberyards[940]}), .top({trees[941], lumberyards[941]}), .top_right({trees[942], lumberyards[942]}), .left({trees[990], lumberyards[990]}), .right({trees[992], lumberyards[992]}), .bottom_left({trees[1040], lumberyards[1040]}), .bottom({trees[1041], lumberyards[1041]}), .bottom_right({trees[1042], lumberyards[1042]}), .init(2'b10), .state({trees[991], lumberyards[991]}));
acre acre_19_42 (.clk(clk), .en(en), .top_left({trees[941], lumberyards[941]}), .top({trees[942], lumberyards[942]}), .top_right({trees[943], lumberyards[943]}), .left({trees[991], lumberyards[991]}), .right({trees[993], lumberyards[993]}), .bottom_left({trees[1041], lumberyards[1041]}), .bottom({trees[1042], lumberyards[1042]}), .bottom_right({trees[1043], lumberyards[1043]}), .init(2'b00), .state({trees[992], lumberyards[992]}));
acre acre_19_43 (.clk(clk), .en(en), .top_left({trees[942], lumberyards[942]}), .top({trees[943], lumberyards[943]}), .top_right({trees[944], lumberyards[944]}), .left({trees[992], lumberyards[992]}), .right({trees[994], lumberyards[994]}), .bottom_left({trees[1042], lumberyards[1042]}), .bottom({trees[1043], lumberyards[1043]}), .bottom_right({trees[1044], lumberyards[1044]}), .init(2'b01), .state({trees[993], lumberyards[993]}));
acre acre_19_44 (.clk(clk), .en(en), .top_left({trees[943], lumberyards[943]}), .top({trees[944], lumberyards[944]}), .top_right({trees[945], lumberyards[945]}), .left({trees[993], lumberyards[993]}), .right({trees[995], lumberyards[995]}), .bottom_left({trees[1043], lumberyards[1043]}), .bottom({trees[1044], lumberyards[1044]}), .bottom_right({trees[1045], lumberyards[1045]}), .init(2'b01), .state({trees[994], lumberyards[994]}));
acre acre_19_45 (.clk(clk), .en(en), .top_left({trees[944], lumberyards[944]}), .top({trees[945], lumberyards[945]}), .top_right({trees[946], lumberyards[946]}), .left({trees[994], lumberyards[994]}), .right({trees[996], lumberyards[996]}), .bottom_left({trees[1044], lumberyards[1044]}), .bottom({trees[1045], lumberyards[1045]}), .bottom_right({trees[1046], lumberyards[1046]}), .init(2'b01), .state({trees[995], lumberyards[995]}));
acre acre_19_46 (.clk(clk), .en(en), .top_left({trees[945], lumberyards[945]}), .top({trees[946], lumberyards[946]}), .top_right({trees[947], lumberyards[947]}), .left({trees[995], lumberyards[995]}), .right({trees[997], lumberyards[997]}), .bottom_left({trees[1045], lumberyards[1045]}), .bottom({trees[1046], lumberyards[1046]}), .bottom_right({trees[1047], lumberyards[1047]}), .init(2'b01), .state({trees[996], lumberyards[996]}));
acre acre_19_47 (.clk(clk), .en(en), .top_left({trees[946], lumberyards[946]}), .top({trees[947], lumberyards[947]}), .top_right({trees[948], lumberyards[948]}), .left({trees[996], lumberyards[996]}), .right({trees[998], lumberyards[998]}), .bottom_left({trees[1046], lumberyards[1046]}), .bottom({trees[1047], lumberyards[1047]}), .bottom_right({trees[1048], lumberyards[1048]}), .init(2'b00), .state({trees[997], lumberyards[997]}));
acre acre_19_48 (.clk(clk), .en(en), .top_left({trees[947], lumberyards[947]}), .top({trees[948], lumberyards[948]}), .top_right({trees[949], lumberyards[949]}), .left({trees[997], lumberyards[997]}), .right({trees[999], lumberyards[999]}), .bottom_left({trees[1047], lumberyards[1047]}), .bottom({trees[1048], lumberyards[1048]}), .bottom_right({trees[1049], lumberyards[1049]}), .init(2'b00), .state({trees[998], lumberyards[998]}));
acre acre_19_49 (.clk(clk), .en(en), .top_left({trees[948], lumberyards[948]}), .top({trees[949], lumberyards[949]}), .top_right(2'b0), .left({trees[998], lumberyards[998]}), .right(2'b0), .bottom_left({trees[1048], lumberyards[1048]}), .bottom({trees[1049], lumberyards[1049]}), .bottom_right(2'b0), .init(2'b00), .state({trees[999], lumberyards[999]}));
acre acre_20_0 (.clk(clk), .en(en), .top_left(2'b0), .top({trees[950], lumberyards[950]}), .top_right({trees[951], lumberyards[951]}), .left(2'b0), .right({trees[1001], lumberyards[1001]}), .bottom_left(2'b0), .bottom({trees[1050], lumberyards[1050]}), .bottom_right({trees[1051], lumberyards[1051]}), .init(2'b00), .state({trees[1000], lumberyards[1000]}));
acre acre_20_1 (.clk(clk), .en(en), .top_left({trees[950], lumberyards[950]}), .top({trees[951], lumberyards[951]}), .top_right({trees[952], lumberyards[952]}), .left({trees[1000], lumberyards[1000]}), .right({trees[1002], lumberyards[1002]}), .bottom_left({trees[1050], lumberyards[1050]}), .bottom({trees[1051], lumberyards[1051]}), .bottom_right({trees[1052], lumberyards[1052]}), .init(2'b00), .state({trees[1001], lumberyards[1001]}));
acre acre_20_2 (.clk(clk), .en(en), .top_left({trees[951], lumberyards[951]}), .top({trees[952], lumberyards[952]}), .top_right({trees[953], lumberyards[953]}), .left({trees[1001], lumberyards[1001]}), .right({trees[1003], lumberyards[1003]}), .bottom_left({trees[1051], lumberyards[1051]}), .bottom({trees[1052], lumberyards[1052]}), .bottom_right({trees[1053], lumberyards[1053]}), .init(2'b00), .state({trees[1002], lumberyards[1002]}));
acre acre_20_3 (.clk(clk), .en(en), .top_left({trees[952], lumberyards[952]}), .top({trees[953], lumberyards[953]}), .top_right({trees[954], lumberyards[954]}), .left({trees[1002], lumberyards[1002]}), .right({trees[1004], lumberyards[1004]}), .bottom_left({trees[1052], lumberyards[1052]}), .bottom({trees[1053], lumberyards[1053]}), .bottom_right({trees[1054], lumberyards[1054]}), .init(2'b00), .state({trees[1003], lumberyards[1003]}));
acre acre_20_4 (.clk(clk), .en(en), .top_left({trees[953], lumberyards[953]}), .top({trees[954], lumberyards[954]}), .top_right({trees[955], lumberyards[955]}), .left({trees[1003], lumberyards[1003]}), .right({trees[1005], lumberyards[1005]}), .bottom_left({trees[1053], lumberyards[1053]}), .bottom({trees[1054], lumberyards[1054]}), .bottom_right({trees[1055], lumberyards[1055]}), .init(2'b00), .state({trees[1004], lumberyards[1004]}));
acre acre_20_5 (.clk(clk), .en(en), .top_left({trees[954], lumberyards[954]}), .top({trees[955], lumberyards[955]}), .top_right({trees[956], lumberyards[956]}), .left({trees[1004], lumberyards[1004]}), .right({trees[1006], lumberyards[1006]}), .bottom_left({trees[1054], lumberyards[1054]}), .bottom({trees[1055], lumberyards[1055]}), .bottom_right({trees[1056], lumberyards[1056]}), .init(2'b00), .state({trees[1005], lumberyards[1005]}));
acre acre_20_6 (.clk(clk), .en(en), .top_left({trees[955], lumberyards[955]}), .top({trees[956], lumberyards[956]}), .top_right({trees[957], lumberyards[957]}), .left({trees[1005], lumberyards[1005]}), .right({trees[1007], lumberyards[1007]}), .bottom_left({trees[1055], lumberyards[1055]}), .bottom({trees[1056], lumberyards[1056]}), .bottom_right({trees[1057], lumberyards[1057]}), .init(2'b10), .state({trees[1006], lumberyards[1006]}));
acre acre_20_7 (.clk(clk), .en(en), .top_left({trees[956], lumberyards[956]}), .top({trees[957], lumberyards[957]}), .top_right({trees[958], lumberyards[958]}), .left({trees[1006], lumberyards[1006]}), .right({trees[1008], lumberyards[1008]}), .bottom_left({trees[1056], lumberyards[1056]}), .bottom({trees[1057], lumberyards[1057]}), .bottom_right({trees[1058], lumberyards[1058]}), .init(2'b00), .state({trees[1007], lumberyards[1007]}));
acre acre_20_8 (.clk(clk), .en(en), .top_left({trees[957], lumberyards[957]}), .top({trees[958], lumberyards[958]}), .top_right({trees[959], lumberyards[959]}), .left({trees[1007], lumberyards[1007]}), .right({trees[1009], lumberyards[1009]}), .bottom_left({trees[1057], lumberyards[1057]}), .bottom({trees[1058], lumberyards[1058]}), .bottom_right({trees[1059], lumberyards[1059]}), .init(2'b10), .state({trees[1008], lumberyards[1008]}));
acre acre_20_9 (.clk(clk), .en(en), .top_left({trees[958], lumberyards[958]}), .top({trees[959], lumberyards[959]}), .top_right({trees[960], lumberyards[960]}), .left({trees[1008], lumberyards[1008]}), .right({trees[1010], lumberyards[1010]}), .bottom_left({trees[1058], lumberyards[1058]}), .bottom({trees[1059], lumberyards[1059]}), .bottom_right({trees[1060], lumberyards[1060]}), .init(2'b00), .state({trees[1009], lumberyards[1009]}));
acre acre_20_10 (.clk(clk), .en(en), .top_left({trees[959], lumberyards[959]}), .top({trees[960], lumberyards[960]}), .top_right({trees[961], lumberyards[961]}), .left({trees[1009], lumberyards[1009]}), .right({trees[1011], lumberyards[1011]}), .bottom_left({trees[1059], lumberyards[1059]}), .bottom({trees[1060], lumberyards[1060]}), .bottom_right({trees[1061], lumberyards[1061]}), .init(2'b10), .state({trees[1010], lumberyards[1010]}));
acre acre_20_11 (.clk(clk), .en(en), .top_left({trees[960], lumberyards[960]}), .top({trees[961], lumberyards[961]}), .top_right({trees[962], lumberyards[962]}), .left({trees[1010], lumberyards[1010]}), .right({trees[1012], lumberyards[1012]}), .bottom_left({trees[1060], lumberyards[1060]}), .bottom({trees[1061], lumberyards[1061]}), .bottom_right({trees[1062], lumberyards[1062]}), .init(2'b10), .state({trees[1011], lumberyards[1011]}));
acre acre_20_12 (.clk(clk), .en(en), .top_left({trees[961], lumberyards[961]}), .top({trees[962], lumberyards[962]}), .top_right({trees[963], lumberyards[963]}), .left({trees[1011], lumberyards[1011]}), .right({trees[1013], lumberyards[1013]}), .bottom_left({trees[1061], lumberyards[1061]}), .bottom({trees[1062], lumberyards[1062]}), .bottom_right({trees[1063], lumberyards[1063]}), .init(2'b00), .state({trees[1012], lumberyards[1012]}));
acre acre_20_13 (.clk(clk), .en(en), .top_left({trees[962], lumberyards[962]}), .top({trees[963], lumberyards[963]}), .top_right({trees[964], lumberyards[964]}), .left({trees[1012], lumberyards[1012]}), .right({trees[1014], lumberyards[1014]}), .bottom_left({trees[1062], lumberyards[1062]}), .bottom({trees[1063], lumberyards[1063]}), .bottom_right({trees[1064], lumberyards[1064]}), .init(2'b10), .state({trees[1013], lumberyards[1013]}));
acre acre_20_14 (.clk(clk), .en(en), .top_left({trees[963], lumberyards[963]}), .top({trees[964], lumberyards[964]}), .top_right({trees[965], lumberyards[965]}), .left({trees[1013], lumberyards[1013]}), .right({trees[1015], lumberyards[1015]}), .bottom_left({trees[1063], lumberyards[1063]}), .bottom({trees[1064], lumberyards[1064]}), .bottom_right({trees[1065], lumberyards[1065]}), .init(2'b10), .state({trees[1014], lumberyards[1014]}));
acre acre_20_15 (.clk(clk), .en(en), .top_left({trees[964], lumberyards[964]}), .top({trees[965], lumberyards[965]}), .top_right({trees[966], lumberyards[966]}), .left({trees[1014], lumberyards[1014]}), .right({trees[1016], lumberyards[1016]}), .bottom_left({trees[1064], lumberyards[1064]}), .bottom({trees[1065], lumberyards[1065]}), .bottom_right({trees[1066], lumberyards[1066]}), .init(2'b00), .state({trees[1015], lumberyards[1015]}));
acre acre_20_16 (.clk(clk), .en(en), .top_left({trees[965], lumberyards[965]}), .top({trees[966], lumberyards[966]}), .top_right({trees[967], lumberyards[967]}), .left({trees[1015], lumberyards[1015]}), .right({trees[1017], lumberyards[1017]}), .bottom_left({trees[1065], lumberyards[1065]}), .bottom({trees[1066], lumberyards[1066]}), .bottom_right({trees[1067], lumberyards[1067]}), .init(2'b01), .state({trees[1016], lumberyards[1016]}));
acre acre_20_17 (.clk(clk), .en(en), .top_left({trees[966], lumberyards[966]}), .top({trees[967], lumberyards[967]}), .top_right({trees[968], lumberyards[968]}), .left({trees[1016], lumberyards[1016]}), .right({trees[1018], lumberyards[1018]}), .bottom_left({trees[1066], lumberyards[1066]}), .bottom({trees[1067], lumberyards[1067]}), .bottom_right({trees[1068], lumberyards[1068]}), .init(2'b01), .state({trees[1017], lumberyards[1017]}));
acre acre_20_18 (.clk(clk), .en(en), .top_left({trees[967], lumberyards[967]}), .top({trees[968], lumberyards[968]}), .top_right({trees[969], lumberyards[969]}), .left({trees[1017], lumberyards[1017]}), .right({trees[1019], lumberyards[1019]}), .bottom_left({trees[1067], lumberyards[1067]}), .bottom({trees[1068], lumberyards[1068]}), .bottom_right({trees[1069], lumberyards[1069]}), .init(2'b01), .state({trees[1018], lumberyards[1018]}));
acre acre_20_19 (.clk(clk), .en(en), .top_left({trees[968], lumberyards[968]}), .top({trees[969], lumberyards[969]}), .top_right({trees[970], lumberyards[970]}), .left({trees[1018], lumberyards[1018]}), .right({trees[1020], lumberyards[1020]}), .bottom_left({trees[1068], lumberyards[1068]}), .bottom({trees[1069], lumberyards[1069]}), .bottom_right({trees[1070], lumberyards[1070]}), .init(2'b00), .state({trees[1019], lumberyards[1019]}));
acre acre_20_20 (.clk(clk), .en(en), .top_left({trees[969], lumberyards[969]}), .top({trees[970], lumberyards[970]}), .top_right({trees[971], lumberyards[971]}), .left({trees[1019], lumberyards[1019]}), .right({trees[1021], lumberyards[1021]}), .bottom_left({trees[1069], lumberyards[1069]}), .bottom({trees[1070], lumberyards[1070]}), .bottom_right({trees[1071], lumberyards[1071]}), .init(2'b01), .state({trees[1020], lumberyards[1020]}));
acre acre_20_21 (.clk(clk), .en(en), .top_left({trees[970], lumberyards[970]}), .top({trees[971], lumberyards[971]}), .top_right({trees[972], lumberyards[972]}), .left({trees[1020], lumberyards[1020]}), .right({trees[1022], lumberyards[1022]}), .bottom_left({trees[1070], lumberyards[1070]}), .bottom({trees[1071], lumberyards[1071]}), .bottom_right({trees[1072], lumberyards[1072]}), .init(2'b00), .state({trees[1021], lumberyards[1021]}));
acre acre_20_22 (.clk(clk), .en(en), .top_left({trees[971], lumberyards[971]}), .top({trees[972], lumberyards[972]}), .top_right({trees[973], lumberyards[973]}), .left({trees[1021], lumberyards[1021]}), .right({trees[1023], lumberyards[1023]}), .bottom_left({trees[1071], lumberyards[1071]}), .bottom({trees[1072], lumberyards[1072]}), .bottom_right({trees[1073], lumberyards[1073]}), .init(2'b01), .state({trees[1022], lumberyards[1022]}));
acre acre_20_23 (.clk(clk), .en(en), .top_left({trees[972], lumberyards[972]}), .top({trees[973], lumberyards[973]}), .top_right({trees[974], lumberyards[974]}), .left({trees[1022], lumberyards[1022]}), .right({trees[1024], lumberyards[1024]}), .bottom_left({trees[1072], lumberyards[1072]}), .bottom({trees[1073], lumberyards[1073]}), .bottom_right({trees[1074], lumberyards[1074]}), .init(2'b01), .state({trees[1023], lumberyards[1023]}));
acre acre_20_24 (.clk(clk), .en(en), .top_left({trees[973], lumberyards[973]}), .top({trees[974], lumberyards[974]}), .top_right({trees[975], lumberyards[975]}), .left({trees[1023], lumberyards[1023]}), .right({trees[1025], lumberyards[1025]}), .bottom_left({trees[1073], lumberyards[1073]}), .bottom({trees[1074], lumberyards[1074]}), .bottom_right({trees[1075], lumberyards[1075]}), .init(2'b01), .state({trees[1024], lumberyards[1024]}));
acre acre_20_25 (.clk(clk), .en(en), .top_left({trees[974], lumberyards[974]}), .top({trees[975], lumberyards[975]}), .top_right({trees[976], lumberyards[976]}), .left({trees[1024], lumberyards[1024]}), .right({trees[1026], lumberyards[1026]}), .bottom_left({trees[1074], lumberyards[1074]}), .bottom({trees[1075], lumberyards[1075]}), .bottom_right({trees[1076], lumberyards[1076]}), .init(2'b00), .state({trees[1025], lumberyards[1025]}));
acre acre_20_26 (.clk(clk), .en(en), .top_left({trees[975], lumberyards[975]}), .top({trees[976], lumberyards[976]}), .top_right({trees[977], lumberyards[977]}), .left({trees[1025], lumberyards[1025]}), .right({trees[1027], lumberyards[1027]}), .bottom_left({trees[1075], lumberyards[1075]}), .bottom({trees[1076], lumberyards[1076]}), .bottom_right({trees[1077], lumberyards[1077]}), .init(2'b00), .state({trees[1026], lumberyards[1026]}));
acre acre_20_27 (.clk(clk), .en(en), .top_left({trees[976], lumberyards[976]}), .top({trees[977], lumberyards[977]}), .top_right({trees[978], lumberyards[978]}), .left({trees[1026], lumberyards[1026]}), .right({trees[1028], lumberyards[1028]}), .bottom_left({trees[1076], lumberyards[1076]}), .bottom({trees[1077], lumberyards[1077]}), .bottom_right({trees[1078], lumberyards[1078]}), .init(2'b00), .state({trees[1027], lumberyards[1027]}));
acre acre_20_28 (.clk(clk), .en(en), .top_left({trees[977], lumberyards[977]}), .top({trees[978], lumberyards[978]}), .top_right({trees[979], lumberyards[979]}), .left({trees[1027], lumberyards[1027]}), .right({trees[1029], lumberyards[1029]}), .bottom_left({trees[1077], lumberyards[1077]}), .bottom({trees[1078], lumberyards[1078]}), .bottom_right({trees[1079], lumberyards[1079]}), .init(2'b00), .state({trees[1028], lumberyards[1028]}));
acre acre_20_29 (.clk(clk), .en(en), .top_left({trees[978], lumberyards[978]}), .top({trees[979], lumberyards[979]}), .top_right({trees[980], lumberyards[980]}), .left({trees[1028], lumberyards[1028]}), .right({trees[1030], lumberyards[1030]}), .bottom_left({trees[1078], lumberyards[1078]}), .bottom({trees[1079], lumberyards[1079]}), .bottom_right({trees[1080], lumberyards[1080]}), .init(2'b00), .state({trees[1029], lumberyards[1029]}));
acre acre_20_30 (.clk(clk), .en(en), .top_left({trees[979], lumberyards[979]}), .top({trees[980], lumberyards[980]}), .top_right({trees[981], lumberyards[981]}), .left({trees[1029], lumberyards[1029]}), .right({trees[1031], lumberyards[1031]}), .bottom_left({trees[1079], lumberyards[1079]}), .bottom({trees[1080], lumberyards[1080]}), .bottom_right({trees[1081], lumberyards[1081]}), .init(2'b00), .state({trees[1030], lumberyards[1030]}));
acre acre_20_31 (.clk(clk), .en(en), .top_left({trees[980], lumberyards[980]}), .top({trees[981], lumberyards[981]}), .top_right({trees[982], lumberyards[982]}), .left({trees[1030], lumberyards[1030]}), .right({trees[1032], lumberyards[1032]}), .bottom_left({trees[1080], lumberyards[1080]}), .bottom({trees[1081], lumberyards[1081]}), .bottom_right({trees[1082], lumberyards[1082]}), .init(2'b00), .state({trees[1031], lumberyards[1031]}));
acre acre_20_32 (.clk(clk), .en(en), .top_left({trees[981], lumberyards[981]}), .top({trees[982], lumberyards[982]}), .top_right({trees[983], lumberyards[983]}), .left({trees[1031], lumberyards[1031]}), .right({trees[1033], lumberyards[1033]}), .bottom_left({trees[1081], lumberyards[1081]}), .bottom({trees[1082], lumberyards[1082]}), .bottom_right({trees[1083], lumberyards[1083]}), .init(2'b00), .state({trees[1032], lumberyards[1032]}));
acre acre_20_33 (.clk(clk), .en(en), .top_left({trees[982], lumberyards[982]}), .top({trees[983], lumberyards[983]}), .top_right({trees[984], lumberyards[984]}), .left({trees[1032], lumberyards[1032]}), .right({trees[1034], lumberyards[1034]}), .bottom_left({trees[1082], lumberyards[1082]}), .bottom({trees[1083], lumberyards[1083]}), .bottom_right({trees[1084], lumberyards[1084]}), .init(2'b00), .state({trees[1033], lumberyards[1033]}));
acre acre_20_34 (.clk(clk), .en(en), .top_left({trees[983], lumberyards[983]}), .top({trees[984], lumberyards[984]}), .top_right({trees[985], lumberyards[985]}), .left({trees[1033], lumberyards[1033]}), .right({trees[1035], lumberyards[1035]}), .bottom_left({trees[1083], lumberyards[1083]}), .bottom({trees[1084], lumberyards[1084]}), .bottom_right({trees[1085], lumberyards[1085]}), .init(2'b00), .state({trees[1034], lumberyards[1034]}));
acre acre_20_35 (.clk(clk), .en(en), .top_left({trees[984], lumberyards[984]}), .top({trees[985], lumberyards[985]}), .top_right({trees[986], lumberyards[986]}), .left({trees[1034], lumberyards[1034]}), .right({trees[1036], lumberyards[1036]}), .bottom_left({trees[1084], lumberyards[1084]}), .bottom({trees[1085], lumberyards[1085]}), .bottom_right({trees[1086], lumberyards[1086]}), .init(2'b01), .state({trees[1035], lumberyards[1035]}));
acre acre_20_36 (.clk(clk), .en(en), .top_left({trees[985], lumberyards[985]}), .top({trees[986], lumberyards[986]}), .top_right({trees[987], lumberyards[987]}), .left({trees[1035], lumberyards[1035]}), .right({trees[1037], lumberyards[1037]}), .bottom_left({trees[1085], lumberyards[1085]}), .bottom({trees[1086], lumberyards[1086]}), .bottom_right({trees[1087], lumberyards[1087]}), .init(2'b00), .state({trees[1036], lumberyards[1036]}));
acre acre_20_37 (.clk(clk), .en(en), .top_left({trees[986], lumberyards[986]}), .top({trees[987], lumberyards[987]}), .top_right({trees[988], lumberyards[988]}), .left({trees[1036], lumberyards[1036]}), .right({trees[1038], lumberyards[1038]}), .bottom_left({trees[1086], lumberyards[1086]}), .bottom({trees[1087], lumberyards[1087]}), .bottom_right({trees[1088], lumberyards[1088]}), .init(2'b00), .state({trees[1037], lumberyards[1037]}));
acre acre_20_38 (.clk(clk), .en(en), .top_left({trees[987], lumberyards[987]}), .top({trees[988], lumberyards[988]}), .top_right({trees[989], lumberyards[989]}), .left({trees[1037], lumberyards[1037]}), .right({trees[1039], lumberyards[1039]}), .bottom_left({trees[1087], lumberyards[1087]}), .bottom({trees[1088], lumberyards[1088]}), .bottom_right({trees[1089], lumberyards[1089]}), .init(2'b00), .state({trees[1038], lumberyards[1038]}));
acre acre_20_39 (.clk(clk), .en(en), .top_left({trees[988], lumberyards[988]}), .top({trees[989], lumberyards[989]}), .top_right({trees[990], lumberyards[990]}), .left({trees[1038], lumberyards[1038]}), .right({trees[1040], lumberyards[1040]}), .bottom_left({trees[1088], lumberyards[1088]}), .bottom({trees[1089], lumberyards[1089]}), .bottom_right({trees[1090], lumberyards[1090]}), .init(2'b10), .state({trees[1039], lumberyards[1039]}));
acre acre_20_40 (.clk(clk), .en(en), .top_left({trees[989], lumberyards[989]}), .top({trees[990], lumberyards[990]}), .top_right({trees[991], lumberyards[991]}), .left({trees[1039], lumberyards[1039]}), .right({trees[1041], lumberyards[1041]}), .bottom_left({trees[1089], lumberyards[1089]}), .bottom({trees[1090], lumberyards[1090]}), .bottom_right({trees[1091], lumberyards[1091]}), .init(2'b10), .state({trees[1040], lumberyards[1040]}));
acre acre_20_41 (.clk(clk), .en(en), .top_left({trees[990], lumberyards[990]}), .top({trees[991], lumberyards[991]}), .top_right({trees[992], lumberyards[992]}), .left({trees[1040], lumberyards[1040]}), .right({trees[1042], lumberyards[1042]}), .bottom_left({trees[1090], lumberyards[1090]}), .bottom({trees[1091], lumberyards[1091]}), .bottom_right({trees[1092], lumberyards[1092]}), .init(2'b10), .state({trees[1041], lumberyards[1041]}));
acre acre_20_42 (.clk(clk), .en(en), .top_left({trees[991], lumberyards[991]}), .top({trees[992], lumberyards[992]}), .top_right({trees[993], lumberyards[993]}), .left({trees[1041], lumberyards[1041]}), .right({trees[1043], lumberyards[1043]}), .bottom_left({trees[1091], lumberyards[1091]}), .bottom({trees[1092], lumberyards[1092]}), .bottom_right({trees[1093], lumberyards[1093]}), .init(2'b00), .state({trees[1042], lumberyards[1042]}));
acre acre_20_43 (.clk(clk), .en(en), .top_left({trees[992], lumberyards[992]}), .top({trees[993], lumberyards[993]}), .top_right({trees[994], lumberyards[994]}), .left({trees[1042], lumberyards[1042]}), .right({trees[1044], lumberyards[1044]}), .bottom_left({trees[1092], lumberyards[1092]}), .bottom({trees[1093], lumberyards[1093]}), .bottom_right({trees[1094], lumberyards[1094]}), .init(2'b00), .state({trees[1043], lumberyards[1043]}));
acre acre_20_44 (.clk(clk), .en(en), .top_left({trees[993], lumberyards[993]}), .top({trees[994], lumberyards[994]}), .top_right({trees[995], lumberyards[995]}), .left({trees[1043], lumberyards[1043]}), .right({trees[1045], lumberyards[1045]}), .bottom_left({trees[1093], lumberyards[1093]}), .bottom({trees[1094], lumberyards[1094]}), .bottom_right({trees[1095], lumberyards[1095]}), .init(2'b00), .state({trees[1044], lumberyards[1044]}));
acre acre_20_45 (.clk(clk), .en(en), .top_left({trees[994], lumberyards[994]}), .top({trees[995], lumberyards[995]}), .top_right({trees[996], lumberyards[996]}), .left({trees[1044], lumberyards[1044]}), .right({trees[1046], lumberyards[1046]}), .bottom_left({trees[1094], lumberyards[1094]}), .bottom({trees[1095], lumberyards[1095]}), .bottom_right({trees[1096], lumberyards[1096]}), .init(2'b01), .state({trees[1045], lumberyards[1045]}));
acre acre_20_46 (.clk(clk), .en(en), .top_left({trees[995], lumberyards[995]}), .top({trees[996], lumberyards[996]}), .top_right({trees[997], lumberyards[997]}), .left({trees[1045], lumberyards[1045]}), .right({trees[1047], lumberyards[1047]}), .bottom_left({trees[1095], lumberyards[1095]}), .bottom({trees[1096], lumberyards[1096]}), .bottom_right({trees[1097], lumberyards[1097]}), .init(2'b01), .state({trees[1046], lumberyards[1046]}));
acre acre_20_47 (.clk(clk), .en(en), .top_left({trees[996], lumberyards[996]}), .top({trees[997], lumberyards[997]}), .top_right({trees[998], lumberyards[998]}), .left({trees[1046], lumberyards[1046]}), .right({trees[1048], lumberyards[1048]}), .bottom_left({trees[1096], lumberyards[1096]}), .bottom({trees[1097], lumberyards[1097]}), .bottom_right({trees[1098], lumberyards[1098]}), .init(2'b01), .state({trees[1047], lumberyards[1047]}));
acre acre_20_48 (.clk(clk), .en(en), .top_left({trees[997], lumberyards[997]}), .top({trees[998], lumberyards[998]}), .top_right({trees[999], lumberyards[999]}), .left({trees[1047], lumberyards[1047]}), .right({trees[1049], lumberyards[1049]}), .bottom_left({trees[1097], lumberyards[1097]}), .bottom({trees[1098], lumberyards[1098]}), .bottom_right({trees[1099], lumberyards[1099]}), .init(2'b00), .state({trees[1048], lumberyards[1048]}));
acre acre_20_49 (.clk(clk), .en(en), .top_left({trees[998], lumberyards[998]}), .top({trees[999], lumberyards[999]}), .top_right(2'b0), .left({trees[1048], lumberyards[1048]}), .right(2'b0), .bottom_left({trees[1098], lumberyards[1098]}), .bottom({trees[1099], lumberyards[1099]}), .bottom_right(2'b0), .init(2'b00), .state({trees[1049], lumberyards[1049]}));
acre acre_21_0 (.clk(clk), .en(en), .top_left(2'b0), .top({trees[1000], lumberyards[1000]}), .top_right({trees[1001], lumberyards[1001]}), .left(2'b0), .right({trees[1051], lumberyards[1051]}), .bottom_left(2'b0), .bottom({trees[1100], lumberyards[1100]}), .bottom_right({trees[1101], lumberyards[1101]}), .init(2'b00), .state({trees[1050], lumberyards[1050]}));
acre acre_21_1 (.clk(clk), .en(en), .top_left({trees[1000], lumberyards[1000]}), .top({trees[1001], lumberyards[1001]}), .top_right({trees[1002], lumberyards[1002]}), .left({trees[1050], lumberyards[1050]}), .right({trees[1052], lumberyards[1052]}), .bottom_left({trees[1100], lumberyards[1100]}), .bottom({trees[1101], lumberyards[1101]}), .bottom_right({trees[1102], lumberyards[1102]}), .init(2'b01), .state({trees[1051], lumberyards[1051]}));
acre acre_21_2 (.clk(clk), .en(en), .top_left({trees[1001], lumberyards[1001]}), .top({trees[1002], lumberyards[1002]}), .top_right({trees[1003], lumberyards[1003]}), .left({trees[1051], lumberyards[1051]}), .right({trees[1053], lumberyards[1053]}), .bottom_left({trees[1101], lumberyards[1101]}), .bottom({trees[1102], lumberyards[1102]}), .bottom_right({trees[1103], lumberyards[1103]}), .init(2'b01), .state({trees[1052], lumberyards[1052]}));
acre acre_21_3 (.clk(clk), .en(en), .top_left({trees[1002], lumberyards[1002]}), .top({trees[1003], lumberyards[1003]}), .top_right({trees[1004], lumberyards[1004]}), .left({trees[1052], lumberyards[1052]}), .right({trees[1054], lumberyards[1054]}), .bottom_left({trees[1102], lumberyards[1102]}), .bottom({trees[1103], lumberyards[1103]}), .bottom_right({trees[1104], lumberyards[1104]}), .init(2'b00), .state({trees[1053], lumberyards[1053]}));
acre acre_21_4 (.clk(clk), .en(en), .top_left({trees[1003], lumberyards[1003]}), .top({trees[1004], lumberyards[1004]}), .top_right({trees[1005], lumberyards[1005]}), .left({trees[1053], lumberyards[1053]}), .right({trees[1055], lumberyards[1055]}), .bottom_left({trees[1103], lumberyards[1103]}), .bottom({trees[1104], lumberyards[1104]}), .bottom_right({trees[1105], lumberyards[1105]}), .init(2'b10), .state({trees[1054], lumberyards[1054]}));
acre acre_21_5 (.clk(clk), .en(en), .top_left({trees[1004], lumberyards[1004]}), .top({trees[1005], lumberyards[1005]}), .top_right({trees[1006], lumberyards[1006]}), .left({trees[1054], lumberyards[1054]}), .right({trees[1056], lumberyards[1056]}), .bottom_left({trees[1104], lumberyards[1104]}), .bottom({trees[1105], lumberyards[1105]}), .bottom_right({trees[1106], lumberyards[1106]}), .init(2'b00), .state({trees[1055], lumberyards[1055]}));
acre acre_21_6 (.clk(clk), .en(en), .top_left({trees[1005], lumberyards[1005]}), .top({trees[1006], lumberyards[1006]}), .top_right({trees[1007], lumberyards[1007]}), .left({trees[1055], lumberyards[1055]}), .right({trees[1057], lumberyards[1057]}), .bottom_left({trees[1105], lumberyards[1105]}), .bottom({trees[1106], lumberyards[1106]}), .bottom_right({trees[1107], lumberyards[1107]}), .init(2'b00), .state({trees[1056], lumberyards[1056]}));
acre acre_21_7 (.clk(clk), .en(en), .top_left({trees[1006], lumberyards[1006]}), .top({trees[1007], lumberyards[1007]}), .top_right({trees[1008], lumberyards[1008]}), .left({trees[1056], lumberyards[1056]}), .right({trees[1058], lumberyards[1058]}), .bottom_left({trees[1106], lumberyards[1106]}), .bottom({trees[1107], lumberyards[1107]}), .bottom_right({trees[1108], lumberyards[1108]}), .init(2'b00), .state({trees[1057], lumberyards[1057]}));
acre acre_21_8 (.clk(clk), .en(en), .top_left({trees[1007], lumberyards[1007]}), .top({trees[1008], lumberyards[1008]}), .top_right({trees[1009], lumberyards[1009]}), .left({trees[1057], lumberyards[1057]}), .right({trees[1059], lumberyards[1059]}), .bottom_left({trees[1107], lumberyards[1107]}), .bottom({trees[1108], lumberyards[1108]}), .bottom_right({trees[1109], lumberyards[1109]}), .init(2'b01), .state({trees[1058], lumberyards[1058]}));
acre acre_21_9 (.clk(clk), .en(en), .top_left({trees[1008], lumberyards[1008]}), .top({trees[1009], lumberyards[1009]}), .top_right({trees[1010], lumberyards[1010]}), .left({trees[1058], lumberyards[1058]}), .right({trees[1060], lumberyards[1060]}), .bottom_left({trees[1108], lumberyards[1108]}), .bottom({trees[1109], lumberyards[1109]}), .bottom_right({trees[1110], lumberyards[1110]}), .init(2'b10), .state({trees[1059], lumberyards[1059]}));
acre acre_21_10 (.clk(clk), .en(en), .top_left({trees[1009], lumberyards[1009]}), .top({trees[1010], lumberyards[1010]}), .top_right({trees[1011], lumberyards[1011]}), .left({trees[1059], lumberyards[1059]}), .right({trees[1061], lumberyards[1061]}), .bottom_left({trees[1109], lumberyards[1109]}), .bottom({trees[1110], lumberyards[1110]}), .bottom_right({trees[1111], lumberyards[1111]}), .init(2'b00), .state({trees[1060], lumberyards[1060]}));
acre acre_21_11 (.clk(clk), .en(en), .top_left({trees[1010], lumberyards[1010]}), .top({trees[1011], lumberyards[1011]}), .top_right({trees[1012], lumberyards[1012]}), .left({trees[1060], lumberyards[1060]}), .right({trees[1062], lumberyards[1062]}), .bottom_left({trees[1110], lumberyards[1110]}), .bottom({trees[1111], lumberyards[1111]}), .bottom_right({trees[1112], lumberyards[1112]}), .init(2'b00), .state({trees[1061], lumberyards[1061]}));
acre acre_21_12 (.clk(clk), .en(en), .top_left({trees[1011], lumberyards[1011]}), .top({trees[1012], lumberyards[1012]}), .top_right({trees[1013], lumberyards[1013]}), .left({trees[1061], lumberyards[1061]}), .right({trees[1063], lumberyards[1063]}), .bottom_left({trees[1111], lumberyards[1111]}), .bottom({trees[1112], lumberyards[1112]}), .bottom_right({trees[1113], lumberyards[1113]}), .init(2'b01), .state({trees[1062], lumberyards[1062]}));
acre acre_21_13 (.clk(clk), .en(en), .top_left({trees[1012], lumberyards[1012]}), .top({trees[1013], lumberyards[1013]}), .top_right({trees[1014], lumberyards[1014]}), .left({trees[1062], lumberyards[1062]}), .right({trees[1064], lumberyards[1064]}), .bottom_left({trees[1112], lumberyards[1112]}), .bottom({trees[1113], lumberyards[1113]}), .bottom_right({trees[1114], lumberyards[1114]}), .init(2'b00), .state({trees[1063], lumberyards[1063]}));
acre acre_21_14 (.clk(clk), .en(en), .top_left({trees[1013], lumberyards[1013]}), .top({trees[1014], lumberyards[1014]}), .top_right({trees[1015], lumberyards[1015]}), .left({trees[1063], lumberyards[1063]}), .right({trees[1065], lumberyards[1065]}), .bottom_left({trees[1113], lumberyards[1113]}), .bottom({trees[1114], lumberyards[1114]}), .bottom_right({trees[1115], lumberyards[1115]}), .init(2'b00), .state({trees[1064], lumberyards[1064]}));
acre acre_21_15 (.clk(clk), .en(en), .top_left({trees[1014], lumberyards[1014]}), .top({trees[1015], lumberyards[1015]}), .top_right({trees[1016], lumberyards[1016]}), .left({trees[1064], lumberyards[1064]}), .right({trees[1066], lumberyards[1066]}), .bottom_left({trees[1114], lumberyards[1114]}), .bottom({trees[1115], lumberyards[1115]}), .bottom_right({trees[1116], lumberyards[1116]}), .init(2'b00), .state({trees[1065], lumberyards[1065]}));
acre acre_21_16 (.clk(clk), .en(en), .top_left({trees[1015], lumberyards[1015]}), .top({trees[1016], lumberyards[1016]}), .top_right({trees[1017], lumberyards[1017]}), .left({trees[1065], lumberyards[1065]}), .right({trees[1067], lumberyards[1067]}), .bottom_left({trees[1115], lumberyards[1115]}), .bottom({trees[1116], lumberyards[1116]}), .bottom_right({trees[1117], lumberyards[1117]}), .init(2'b00), .state({trees[1066], lumberyards[1066]}));
acre acre_21_17 (.clk(clk), .en(en), .top_left({trees[1016], lumberyards[1016]}), .top({trees[1017], lumberyards[1017]}), .top_right({trees[1018], lumberyards[1018]}), .left({trees[1066], lumberyards[1066]}), .right({trees[1068], lumberyards[1068]}), .bottom_left({trees[1116], lumberyards[1116]}), .bottom({trees[1117], lumberyards[1117]}), .bottom_right({trees[1118], lumberyards[1118]}), .init(2'b10), .state({trees[1067], lumberyards[1067]}));
acre acre_21_18 (.clk(clk), .en(en), .top_left({trees[1017], lumberyards[1017]}), .top({trees[1018], lumberyards[1018]}), .top_right({trees[1019], lumberyards[1019]}), .left({trees[1067], lumberyards[1067]}), .right({trees[1069], lumberyards[1069]}), .bottom_left({trees[1117], lumberyards[1117]}), .bottom({trees[1118], lumberyards[1118]}), .bottom_right({trees[1119], lumberyards[1119]}), .init(2'b00), .state({trees[1068], lumberyards[1068]}));
acre acre_21_19 (.clk(clk), .en(en), .top_left({trees[1018], lumberyards[1018]}), .top({trees[1019], lumberyards[1019]}), .top_right({trees[1020], lumberyards[1020]}), .left({trees[1068], lumberyards[1068]}), .right({trees[1070], lumberyards[1070]}), .bottom_left({trees[1118], lumberyards[1118]}), .bottom({trees[1119], lumberyards[1119]}), .bottom_right({trees[1120], lumberyards[1120]}), .init(2'b01), .state({trees[1069], lumberyards[1069]}));
acre acre_21_20 (.clk(clk), .en(en), .top_left({trees[1019], lumberyards[1019]}), .top({trees[1020], lumberyards[1020]}), .top_right({trees[1021], lumberyards[1021]}), .left({trees[1069], lumberyards[1069]}), .right({trees[1071], lumberyards[1071]}), .bottom_left({trees[1119], lumberyards[1119]}), .bottom({trees[1120], lumberyards[1120]}), .bottom_right({trees[1121], lumberyards[1121]}), .init(2'b00), .state({trees[1070], lumberyards[1070]}));
acre acre_21_21 (.clk(clk), .en(en), .top_left({trees[1020], lumberyards[1020]}), .top({trees[1021], lumberyards[1021]}), .top_right({trees[1022], lumberyards[1022]}), .left({trees[1070], lumberyards[1070]}), .right({trees[1072], lumberyards[1072]}), .bottom_left({trees[1120], lumberyards[1120]}), .bottom({trees[1121], lumberyards[1121]}), .bottom_right({trees[1122], lumberyards[1122]}), .init(2'b00), .state({trees[1071], lumberyards[1071]}));
acre acre_21_22 (.clk(clk), .en(en), .top_left({trees[1021], lumberyards[1021]}), .top({trees[1022], lumberyards[1022]}), .top_right({trees[1023], lumberyards[1023]}), .left({trees[1071], lumberyards[1071]}), .right({trees[1073], lumberyards[1073]}), .bottom_left({trees[1121], lumberyards[1121]}), .bottom({trees[1122], lumberyards[1122]}), .bottom_right({trees[1123], lumberyards[1123]}), .init(2'b00), .state({trees[1072], lumberyards[1072]}));
acre acre_21_23 (.clk(clk), .en(en), .top_left({trees[1022], lumberyards[1022]}), .top({trees[1023], lumberyards[1023]}), .top_right({trees[1024], lumberyards[1024]}), .left({trees[1072], lumberyards[1072]}), .right({trees[1074], lumberyards[1074]}), .bottom_left({trees[1122], lumberyards[1122]}), .bottom({trees[1123], lumberyards[1123]}), .bottom_right({trees[1124], lumberyards[1124]}), .init(2'b01), .state({trees[1073], lumberyards[1073]}));
acre acre_21_24 (.clk(clk), .en(en), .top_left({trees[1023], lumberyards[1023]}), .top({trees[1024], lumberyards[1024]}), .top_right({trees[1025], lumberyards[1025]}), .left({trees[1073], lumberyards[1073]}), .right({trees[1075], lumberyards[1075]}), .bottom_left({trees[1123], lumberyards[1123]}), .bottom({trees[1124], lumberyards[1124]}), .bottom_right({trees[1125], lumberyards[1125]}), .init(2'b00), .state({trees[1074], lumberyards[1074]}));
acre acre_21_25 (.clk(clk), .en(en), .top_left({trees[1024], lumberyards[1024]}), .top({trees[1025], lumberyards[1025]}), .top_right({trees[1026], lumberyards[1026]}), .left({trees[1074], lumberyards[1074]}), .right({trees[1076], lumberyards[1076]}), .bottom_left({trees[1124], lumberyards[1124]}), .bottom({trees[1125], lumberyards[1125]}), .bottom_right({trees[1126], lumberyards[1126]}), .init(2'b00), .state({trees[1075], lumberyards[1075]}));
acre acre_21_26 (.clk(clk), .en(en), .top_left({trees[1025], lumberyards[1025]}), .top({trees[1026], lumberyards[1026]}), .top_right({trees[1027], lumberyards[1027]}), .left({trees[1075], lumberyards[1075]}), .right({trees[1077], lumberyards[1077]}), .bottom_left({trees[1125], lumberyards[1125]}), .bottom({trees[1126], lumberyards[1126]}), .bottom_right({trees[1127], lumberyards[1127]}), .init(2'b00), .state({trees[1076], lumberyards[1076]}));
acre acre_21_27 (.clk(clk), .en(en), .top_left({trees[1026], lumberyards[1026]}), .top({trees[1027], lumberyards[1027]}), .top_right({trees[1028], lumberyards[1028]}), .left({trees[1076], lumberyards[1076]}), .right({trees[1078], lumberyards[1078]}), .bottom_left({trees[1126], lumberyards[1126]}), .bottom({trees[1127], lumberyards[1127]}), .bottom_right({trees[1128], lumberyards[1128]}), .init(2'b01), .state({trees[1077], lumberyards[1077]}));
acre acre_21_28 (.clk(clk), .en(en), .top_left({trees[1027], lumberyards[1027]}), .top({trees[1028], lumberyards[1028]}), .top_right({trees[1029], lumberyards[1029]}), .left({trees[1077], lumberyards[1077]}), .right({trees[1079], lumberyards[1079]}), .bottom_left({trees[1127], lumberyards[1127]}), .bottom({trees[1128], lumberyards[1128]}), .bottom_right({trees[1129], lumberyards[1129]}), .init(2'b10), .state({trees[1078], lumberyards[1078]}));
acre acre_21_29 (.clk(clk), .en(en), .top_left({trees[1028], lumberyards[1028]}), .top({trees[1029], lumberyards[1029]}), .top_right({trees[1030], lumberyards[1030]}), .left({trees[1078], lumberyards[1078]}), .right({trees[1080], lumberyards[1080]}), .bottom_left({trees[1128], lumberyards[1128]}), .bottom({trees[1129], lumberyards[1129]}), .bottom_right({trees[1130], lumberyards[1130]}), .init(2'b00), .state({trees[1079], lumberyards[1079]}));
acre acre_21_30 (.clk(clk), .en(en), .top_left({trees[1029], lumberyards[1029]}), .top({trees[1030], lumberyards[1030]}), .top_right({trees[1031], lumberyards[1031]}), .left({trees[1079], lumberyards[1079]}), .right({trees[1081], lumberyards[1081]}), .bottom_left({trees[1129], lumberyards[1129]}), .bottom({trees[1130], lumberyards[1130]}), .bottom_right({trees[1131], lumberyards[1131]}), .init(2'b01), .state({trees[1080], lumberyards[1080]}));
acre acre_21_31 (.clk(clk), .en(en), .top_left({trees[1030], lumberyards[1030]}), .top({trees[1031], lumberyards[1031]}), .top_right({trees[1032], lumberyards[1032]}), .left({trees[1080], lumberyards[1080]}), .right({trees[1082], lumberyards[1082]}), .bottom_left({trees[1130], lumberyards[1130]}), .bottom({trees[1131], lumberyards[1131]}), .bottom_right({trees[1132], lumberyards[1132]}), .init(2'b01), .state({trees[1081], lumberyards[1081]}));
acre acre_21_32 (.clk(clk), .en(en), .top_left({trees[1031], lumberyards[1031]}), .top({trees[1032], lumberyards[1032]}), .top_right({trees[1033], lumberyards[1033]}), .left({trees[1081], lumberyards[1081]}), .right({trees[1083], lumberyards[1083]}), .bottom_left({trees[1131], lumberyards[1131]}), .bottom({trees[1132], lumberyards[1132]}), .bottom_right({trees[1133], lumberyards[1133]}), .init(2'b00), .state({trees[1082], lumberyards[1082]}));
acre acre_21_33 (.clk(clk), .en(en), .top_left({trees[1032], lumberyards[1032]}), .top({trees[1033], lumberyards[1033]}), .top_right({trees[1034], lumberyards[1034]}), .left({trees[1082], lumberyards[1082]}), .right({trees[1084], lumberyards[1084]}), .bottom_left({trees[1132], lumberyards[1132]}), .bottom({trees[1133], lumberyards[1133]}), .bottom_right({trees[1134], lumberyards[1134]}), .init(2'b10), .state({trees[1083], lumberyards[1083]}));
acre acre_21_34 (.clk(clk), .en(en), .top_left({trees[1033], lumberyards[1033]}), .top({trees[1034], lumberyards[1034]}), .top_right({trees[1035], lumberyards[1035]}), .left({trees[1083], lumberyards[1083]}), .right({trees[1085], lumberyards[1085]}), .bottom_left({trees[1133], lumberyards[1133]}), .bottom({trees[1134], lumberyards[1134]}), .bottom_right({trees[1135], lumberyards[1135]}), .init(2'b01), .state({trees[1084], lumberyards[1084]}));
acre acre_21_35 (.clk(clk), .en(en), .top_left({trees[1034], lumberyards[1034]}), .top({trees[1035], lumberyards[1035]}), .top_right({trees[1036], lumberyards[1036]}), .left({trees[1084], lumberyards[1084]}), .right({trees[1086], lumberyards[1086]}), .bottom_left({trees[1134], lumberyards[1134]}), .bottom({trees[1135], lumberyards[1135]}), .bottom_right({trees[1136], lumberyards[1136]}), .init(2'b00), .state({trees[1085], lumberyards[1085]}));
acre acre_21_36 (.clk(clk), .en(en), .top_left({trees[1035], lumberyards[1035]}), .top({trees[1036], lumberyards[1036]}), .top_right({trees[1037], lumberyards[1037]}), .left({trees[1085], lumberyards[1085]}), .right({trees[1087], lumberyards[1087]}), .bottom_left({trees[1135], lumberyards[1135]}), .bottom({trees[1136], lumberyards[1136]}), .bottom_right({trees[1137], lumberyards[1137]}), .init(2'b10), .state({trees[1086], lumberyards[1086]}));
acre acre_21_37 (.clk(clk), .en(en), .top_left({trees[1036], lumberyards[1036]}), .top({trees[1037], lumberyards[1037]}), .top_right({trees[1038], lumberyards[1038]}), .left({trees[1086], lumberyards[1086]}), .right({trees[1088], lumberyards[1088]}), .bottom_left({trees[1136], lumberyards[1136]}), .bottom({trees[1137], lumberyards[1137]}), .bottom_right({trees[1138], lumberyards[1138]}), .init(2'b10), .state({trees[1087], lumberyards[1087]}));
acre acre_21_38 (.clk(clk), .en(en), .top_left({trees[1037], lumberyards[1037]}), .top({trees[1038], lumberyards[1038]}), .top_right({trees[1039], lumberyards[1039]}), .left({trees[1087], lumberyards[1087]}), .right({trees[1089], lumberyards[1089]}), .bottom_left({trees[1137], lumberyards[1137]}), .bottom({trees[1138], lumberyards[1138]}), .bottom_right({trees[1139], lumberyards[1139]}), .init(2'b00), .state({trees[1088], lumberyards[1088]}));
acre acre_21_39 (.clk(clk), .en(en), .top_left({trees[1038], lumberyards[1038]}), .top({trees[1039], lumberyards[1039]}), .top_right({trees[1040], lumberyards[1040]}), .left({trees[1088], lumberyards[1088]}), .right({trees[1090], lumberyards[1090]}), .bottom_left({trees[1138], lumberyards[1138]}), .bottom({trees[1139], lumberyards[1139]}), .bottom_right({trees[1140], lumberyards[1140]}), .init(2'b00), .state({trees[1089], lumberyards[1089]}));
acre acre_21_40 (.clk(clk), .en(en), .top_left({trees[1039], lumberyards[1039]}), .top({trees[1040], lumberyards[1040]}), .top_right({trees[1041], lumberyards[1041]}), .left({trees[1089], lumberyards[1089]}), .right({trees[1091], lumberyards[1091]}), .bottom_left({trees[1139], lumberyards[1139]}), .bottom({trees[1140], lumberyards[1140]}), .bottom_right({trees[1141], lumberyards[1141]}), .init(2'b01), .state({trees[1090], lumberyards[1090]}));
acre acre_21_41 (.clk(clk), .en(en), .top_left({trees[1040], lumberyards[1040]}), .top({trees[1041], lumberyards[1041]}), .top_right({trees[1042], lumberyards[1042]}), .left({trees[1090], lumberyards[1090]}), .right({trees[1092], lumberyards[1092]}), .bottom_left({trees[1140], lumberyards[1140]}), .bottom({trees[1141], lumberyards[1141]}), .bottom_right({trees[1142], lumberyards[1142]}), .init(2'b00), .state({trees[1091], lumberyards[1091]}));
acre acre_21_42 (.clk(clk), .en(en), .top_left({trees[1041], lumberyards[1041]}), .top({trees[1042], lumberyards[1042]}), .top_right({trees[1043], lumberyards[1043]}), .left({trees[1091], lumberyards[1091]}), .right({trees[1093], lumberyards[1093]}), .bottom_left({trees[1141], lumberyards[1141]}), .bottom({trees[1142], lumberyards[1142]}), .bottom_right({trees[1143], lumberyards[1143]}), .init(2'b10), .state({trees[1092], lumberyards[1092]}));
acre acre_21_43 (.clk(clk), .en(en), .top_left({trees[1042], lumberyards[1042]}), .top({trees[1043], lumberyards[1043]}), .top_right({trees[1044], lumberyards[1044]}), .left({trees[1092], lumberyards[1092]}), .right({trees[1094], lumberyards[1094]}), .bottom_left({trees[1142], lumberyards[1142]}), .bottom({trees[1143], lumberyards[1143]}), .bottom_right({trees[1144], lumberyards[1144]}), .init(2'b00), .state({trees[1093], lumberyards[1093]}));
acre acre_21_44 (.clk(clk), .en(en), .top_left({trees[1043], lumberyards[1043]}), .top({trees[1044], lumberyards[1044]}), .top_right({trees[1045], lumberyards[1045]}), .left({trees[1093], lumberyards[1093]}), .right({trees[1095], lumberyards[1095]}), .bottom_left({trees[1143], lumberyards[1143]}), .bottom({trees[1144], lumberyards[1144]}), .bottom_right({trees[1145], lumberyards[1145]}), .init(2'b00), .state({trees[1094], lumberyards[1094]}));
acre acre_21_45 (.clk(clk), .en(en), .top_left({trees[1044], lumberyards[1044]}), .top({trees[1045], lumberyards[1045]}), .top_right({trees[1046], lumberyards[1046]}), .left({trees[1094], lumberyards[1094]}), .right({trees[1096], lumberyards[1096]}), .bottom_left({trees[1144], lumberyards[1144]}), .bottom({trees[1145], lumberyards[1145]}), .bottom_right({trees[1146], lumberyards[1146]}), .init(2'b10), .state({trees[1095], lumberyards[1095]}));
acre acre_21_46 (.clk(clk), .en(en), .top_left({trees[1045], lumberyards[1045]}), .top({trees[1046], lumberyards[1046]}), .top_right({trees[1047], lumberyards[1047]}), .left({trees[1095], lumberyards[1095]}), .right({trees[1097], lumberyards[1097]}), .bottom_left({trees[1145], lumberyards[1145]}), .bottom({trees[1146], lumberyards[1146]}), .bottom_right({trees[1147], lumberyards[1147]}), .init(2'b00), .state({trees[1096], lumberyards[1096]}));
acre acre_21_47 (.clk(clk), .en(en), .top_left({trees[1046], lumberyards[1046]}), .top({trees[1047], lumberyards[1047]}), .top_right({trees[1048], lumberyards[1048]}), .left({trees[1096], lumberyards[1096]}), .right({trees[1098], lumberyards[1098]}), .bottom_left({trees[1146], lumberyards[1146]}), .bottom({trees[1147], lumberyards[1147]}), .bottom_right({trees[1148], lumberyards[1148]}), .init(2'b10), .state({trees[1097], lumberyards[1097]}));
acre acre_21_48 (.clk(clk), .en(en), .top_left({trees[1047], lumberyards[1047]}), .top({trees[1048], lumberyards[1048]}), .top_right({trees[1049], lumberyards[1049]}), .left({trees[1097], lumberyards[1097]}), .right({trees[1099], lumberyards[1099]}), .bottom_left({trees[1147], lumberyards[1147]}), .bottom({trees[1148], lumberyards[1148]}), .bottom_right({trees[1149], lumberyards[1149]}), .init(2'b01), .state({trees[1098], lumberyards[1098]}));
acre acre_21_49 (.clk(clk), .en(en), .top_left({trees[1048], lumberyards[1048]}), .top({trees[1049], lumberyards[1049]}), .top_right(2'b0), .left({trees[1098], lumberyards[1098]}), .right(2'b0), .bottom_left({trees[1148], lumberyards[1148]}), .bottom({trees[1149], lumberyards[1149]}), .bottom_right(2'b0), .init(2'b00), .state({trees[1099], lumberyards[1099]}));
acre acre_22_0 (.clk(clk), .en(en), .top_left(2'b0), .top({trees[1050], lumberyards[1050]}), .top_right({trees[1051], lumberyards[1051]}), .left(2'b0), .right({trees[1101], lumberyards[1101]}), .bottom_left(2'b0), .bottom({trees[1150], lumberyards[1150]}), .bottom_right({trees[1151], lumberyards[1151]}), .init(2'b10), .state({trees[1100], lumberyards[1100]}));
acre acre_22_1 (.clk(clk), .en(en), .top_left({trees[1050], lumberyards[1050]}), .top({trees[1051], lumberyards[1051]}), .top_right({trees[1052], lumberyards[1052]}), .left({trees[1100], lumberyards[1100]}), .right({trees[1102], lumberyards[1102]}), .bottom_left({trees[1150], lumberyards[1150]}), .bottom({trees[1151], lumberyards[1151]}), .bottom_right({trees[1152], lumberyards[1152]}), .init(2'b10), .state({trees[1101], lumberyards[1101]}));
acre acre_22_2 (.clk(clk), .en(en), .top_left({trees[1051], lumberyards[1051]}), .top({trees[1052], lumberyards[1052]}), .top_right({trees[1053], lumberyards[1053]}), .left({trees[1101], lumberyards[1101]}), .right({trees[1103], lumberyards[1103]}), .bottom_left({trees[1151], lumberyards[1151]}), .bottom({trees[1152], lumberyards[1152]}), .bottom_right({trees[1153], lumberyards[1153]}), .init(2'b00), .state({trees[1102], lumberyards[1102]}));
acre acre_22_3 (.clk(clk), .en(en), .top_left({trees[1052], lumberyards[1052]}), .top({trees[1053], lumberyards[1053]}), .top_right({trees[1054], lumberyards[1054]}), .left({trees[1102], lumberyards[1102]}), .right({trees[1104], lumberyards[1104]}), .bottom_left({trees[1152], lumberyards[1152]}), .bottom({trees[1153], lumberyards[1153]}), .bottom_right({trees[1154], lumberyards[1154]}), .init(2'b00), .state({trees[1103], lumberyards[1103]}));
acre acre_22_4 (.clk(clk), .en(en), .top_left({trees[1053], lumberyards[1053]}), .top({trees[1054], lumberyards[1054]}), .top_right({trees[1055], lumberyards[1055]}), .left({trees[1103], lumberyards[1103]}), .right({trees[1105], lumberyards[1105]}), .bottom_left({trees[1153], lumberyards[1153]}), .bottom({trees[1154], lumberyards[1154]}), .bottom_right({trees[1155], lumberyards[1155]}), .init(2'b00), .state({trees[1104], lumberyards[1104]}));
acre acre_22_5 (.clk(clk), .en(en), .top_left({trees[1054], lumberyards[1054]}), .top({trees[1055], lumberyards[1055]}), .top_right({trees[1056], lumberyards[1056]}), .left({trees[1104], lumberyards[1104]}), .right({trees[1106], lumberyards[1106]}), .bottom_left({trees[1154], lumberyards[1154]}), .bottom({trees[1155], lumberyards[1155]}), .bottom_right({trees[1156], lumberyards[1156]}), .init(2'b00), .state({trees[1105], lumberyards[1105]}));
acre acre_22_6 (.clk(clk), .en(en), .top_left({trees[1055], lumberyards[1055]}), .top({trees[1056], lumberyards[1056]}), .top_right({trees[1057], lumberyards[1057]}), .left({trees[1105], lumberyards[1105]}), .right({trees[1107], lumberyards[1107]}), .bottom_left({trees[1155], lumberyards[1155]}), .bottom({trees[1156], lumberyards[1156]}), .bottom_right({trees[1157], lumberyards[1157]}), .init(2'b01), .state({trees[1106], lumberyards[1106]}));
acre acre_22_7 (.clk(clk), .en(en), .top_left({trees[1056], lumberyards[1056]}), .top({trees[1057], lumberyards[1057]}), .top_right({trees[1058], lumberyards[1058]}), .left({trees[1106], lumberyards[1106]}), .right({trees[1108], lumberyards[1108]}), .bottom_left({trees[1156], lumberyards[1156]}), .bottom({trees[1157], lumberyards[1157]}), .bottom_right({trees[1158], lumberyards[1158]}), .init(2'b10), .state({trees[1107], lumberyards[1107]}));
acre acre_22_8 (.clk(clk), .en(en), .top_left({trees[1057], lumberyards[1057]}), .top({trees[1058], lumberyards[1058]}), .top_right({trees[1059], lumberyards[1059]}), .left({trees[1107], lumberyards[1107]}), .right({trees[1109], lumberyards[1109]}), .bottom_left({trees[1157], lumberyards[1157]}), .bottom({trees[1158], lumberyards[1158]}), .bottom_right({trees[1159], lumberyards[1159]}), .init(2'b01), .state({trees[1108], lumberyards[1108]}));
acre acre_22_9 (.clk(clk), .en(en), .top_left({trees[1058], lumberyards[1058]}), .top({trees[1059], lumberyards[1059]}), .top_right({trees[1060], lumberyards[1060]}), .left({trees[1108], lumberyards[1108]}), .right({trees[1110], lumberyards[1110]}), .bottom_left({trees[1158], lumberyards[1158]}), .bottom({trees[1159], lumberyards[1159]}), .bottom_right({trees[1160], lumberyards[1160]}), .init(2'b10), .state({trees[1109], lumberyards[1109]}));
acre acre_22_10 (.clk(clk), .en(en), .top_left({trees[1059], lumberyards[1059]}), .top({trees[1060], lumberyards[1060]}), .top_right({trees[1061], lumberyards[1061]}), .left({trees[1109], lumberyards[1109]}), .right({trees[1111], lumberyards[1111]}), .bottom_left({trees[1159], lumberyards[1159]}), .bottom({trees[1160], lumberyards[1160]}), .bottom_right({trees[1161], lumberyards[1161]}), .init(2'b00), .state({trees[1110], lumberyards[1110]}));
acre acre_22_11 (.clk(clk), .en(en), .top_left({trees[1060], lumberyards[1060]}), .top({trees[1061], lumberyards[1061]}), .top_right({trees[1062], lumberyards[1062]}), .left({trees[1110], lumberyards[1110]}), .right({trees[1112], lumberyards[1112]}), .bottom_left({trees[1160], lumberyards[1160]}), .bottom({trees[1161], lumberyards[1161]}), .bottom_right({trees[1162], lumberyards[1162]}), .init(2'b01), .state({trees[1111], lumberyards[1111]}));
acre acre_22_12 (.clk(clk), .en(en), .top_left({trees[1061], lumberyards[1061]}), .top({trees[1062], lumberyards[1062]}), .top_right({trees[1063], lumberyards[1063]}), .left({trees[1111], lumberyards[1111]}), .right({trees[1113], lumberyards[1113]}), .bottom_left({trees[1161], lumberyards[1161]}), .bottom({trees[1162], lumberyards[1162]}), .bottom_right({trees[1163], lumberyards[1163]}), .init(2'b10), .state({trees[1112], lumberyards[1112]}));
acre acre_22_13 (.clk(clk), .en(en), .top_left({trees[1062], lumberyards[1062]}), .top({trees[1063], lumberyards[1063]}), .top_right({trees[1064], lumberyards[1064]}), .left({trees[1112], lumberyards[1112]}), .right({trees[1114], lumberyards[1114]}), .bottom_left({trees[1162], lumberyards[1162]}), .bottom({trees[1163], lumberyards[1163]}), .bottom_right({trees[1164], lumberyards[1164]}), .init(2'b10), .state({trees[1113], lumberyards[1113]}));
acre acre_22_14 (.clk(clk), .en(en), .top_left({trees[1063], lumberyards[1063]}), .top({trees[1064], lumberyards[1064]}), .top_right({trees[1065], lumberyards[1065]}), .left({trees[1113], lumberyards[1113]}), .right({trees[1115], lumberyards[1115]}), .bottom_left({trees[1163], lumberyards[1163]}), .bottom({trees[1164], lumberyards[1164]}), .bottom_right({trees[1165], lumberyards[1165]}), .init(2'b10), .state({trees[1114], lumberyards[1114]}));
acre acre_22_15 (.clk(clk), .en(en), .top_left({trees[1064], lumberyards[1064]}), .top({trees[1065], lumberyards[1065]}), .top_right({trees[1066], lumberyards[1066]}), .left({trees[1114], lumberyards[1114]}), .right({trees[1116], lumberyards[1116]}), .bottom_left({trees[1164], lumberyards[1164]}), .bottom({trees[1165], lumberyards[1165]}), .bottom_right({trees[1166], lumberyards[1166]}), .init(2'b00), .state({trees[1115], lumberyards[1115]}));
acre acre_22_16 (.clk(clk), .en(en), .top_left({trees[1065], lumberyards[1065]}), .top({trees[1066], lumberyards[1066]}), .top_right({trees[1067], lumberyards[1067]}), .left({trees[1115], lumberyards[1115]}), .right({trees[1117], lumberyards[1117]}), .bottom_left({trees[1165], lumberyards[1165]}), .bottom({trees[1166], lumberyards[1166]}), .bottom_right({trees[1167], lumberyards[1167]}), .init(2'b10), .state({trees[1116], lumberyards[1116]}));
acre acre_22_17 (.clk(clk), .en(en), .top_left({trees[1066], lumberyards[1066]}), .top({trees[1067], lumberyards[1067]}), .top_right({trees[1068], lumberyards[1068]}), .left({trees[1116], lumberyards[1116]}), .right({trees[1118], lumberyards[1118]}), .bottom_left({trees[1166], lumberyards[1166]}), .bottom({trees[1167], lumberyards[1167]}), .bottom_right({trees[1168], lumberyards[1168]}), .init(2'b00), .state({trees[1117], lumberyards[1117]}));
acre acre_22_18 (.clk(clk), .en(en), .top_left({trees[1067], lumberyards[1067]}), .top({trees[1068], lumberyards[1068]}), .top_right({trees[1069], lumberyards[1069]}), .left({trees[1117], lumberyards[1117]}), .right({trees[1119], lumberyards[1119]}), .bottom_left({trees[1167], lumberyards[1167]}), .bottom({trees[1168], lumberyards[1168]}), .bottom_right({trees[1169], lumberyards[1169]}), .init(2'b00), .state({trees[1118], lumberyards[1118]}));
acre acre_22_19 (.clk(clk), .en(en), .top_left({trees[1068], lumberyards[1068]}), .top({trees[1069], lumberyards[1069]}), .top_right({trees[1070], lumberyards[1070]}), .left({trees[1118], lumberyards[1118]}), .right({trees[1120], lumberyards[1120]}), .bottom_left({trees[1168], lumberyards[1168]}), .bottom({trees[1169], lumberyards[1169]}), .bottom_right({trees[1170], lumberyards[1170]}), .init(2'b00), .state({trees[1119], lumberyards[1119]}));
acre acre_22_20 (.clk(clk), .en(en), .top_left({trees[1069], lumberyards[1069]}), .top({trees[1070], lumberyards[1070]}), .top_right({trees[1071], lumberyards[1071]}), .left({trees[1119], lumberyards[1119]}), .right({trees[1121], lumberyards[1121]}), .bottom_left({trees[1169], lumberyards[1169]}), .bottom({trees[1170], lumberyards[1170]}), .bottom_right({trees[1171], lumberyards[1171]}), .init(2'b10), .state({trees[1120], lumberyards[1120]}));
acre acre_22_21 (.clk(clk), .en(en), .top_left({trees[1070], lumberyards[1070]}), .top({trees[1071], lumberyards[1071]}), .top_right({trees[1072], lumberyards[1072]}), .left({trees[1120], lumberyards[1120]}), .right({trees[1122], lumberyards[1122]}), .bottom_left({trees[1170], lumberyards[1170]}), .bottom({trees[1171], lumberyards[1171]}), .bottom_right({trees[1172], lumberyards[1172]}), .init(2'b10), .state({trees[1121], lumberyards[1121]}));
acre acre_22_22 (.clk(clk), .en(en), .top_left({trees[1071], lumberyards[1071]}), .top({trees[1072], lumberyards[1072]}), .top_right({trees[1073], lumberyards[1073]}), .left({trees[1121], lumberyards[1121]}), .right({trees[1123], lumberyards[1123]}), .bottom_left({trees[1171], lumberyards[1171]}), .bottom({trees[1172], lumberyards[1172]}), .bottom_right({trees[1173], lumberyards[1173]}), .init(2'b00), .state({trees[1122], lumberyards[1122]}));
acre acre_22_23 (.clk(clk), .en(en), .top_left({trees[1072], lumberyards[1072]}), .top({trees[1073], lumberyards[1073]}), .top_right({trees[1074], lumberyards[1074]}), .left({trees[1122], lumberyards[1122]}), .right({trees[1124], lumberyards[1124]}), .bottom_left({trees[1172], lumberyards[1172]}), .bottom({trees[1173], lumberyards[1173]}), .bottom_right({trees[1174], lumberyards[1174]}), .init(2'b00), .state({trees[1123], lumberyards[1123]}));
acre acre_22_24 (.clk(clk), .en(en), .top_left({trees[1073], lumberyards[1073]}), .top({trees[1074], lumberyards[1074]}), .top_right({trees[1075], lumberyards[1075]}), .left({trees[1123], lumberyards[1123]}), .right({trees[1125], lumberyards[1125]}), .bottom_left({trees[1173], lumberyards[1173]}), .bottom({trees[1174], lumberyards[1174]}), .bottom_right({trees[1175], lumberyards[1175]}), .init(2'b10), .state({trees[1124], lumberyards[1124]}));
acre acre_22_25 (.clk(clk), .en(en), .top_left({trees[1074], lumberyards[1074]}), .top({trees[1075], lumberyards[1075]}), .top_right({trees[1076], lumberyards[1076]}), .left({trees[1124], lumberyards[1124]}), .right({trees[1126], lumberyards[1126]}), .bottom_left({trees[1174], lumberyards[1174]}), .bottom({trees[1175], lumberyards[1175]}), .bottom_right({trees[1176], lumberyards[1176]}), .init(2'b00), .state({trees[1125], lumberyards[1125]}));
acre acre_22_26 (.clk(clk), .en(en), .top_left({trees[1075], lumberyards[1075]}), .top({trees[1076], lumberyards[1076]}), .top_right({trees[1077], lumberyards[1077]}), .left({trees[1125], lumberyards[1125]}), .right({trees[1127], lumberyards[1127]}), .bottom_left({trees[1175], lumberyards[1175]}), .bottom({trees[1176], lumberyards[1176]}), .bottom_right({trees[1177], lumberyards[1177]}), .init(2'b01), .state({trees[1126], lumberyards[1126]}));
acre acre_22_27 (.clk(clk), .en(en), .top_left({trees[1076], lumberyards[1076]}), .top({trees[1077], lumberyards[1077]}), .top_right({trees[1078], lumberyards[1078]}), .left({trees[1126], lumberyards[1126]}), .right({trees[1128], lumberyards[1128]}), .bottom_left({trees[1176], lumberyards[1176]}), .bottom({trees[1177], lumberyards[1177]}), .bottom_right({trees[1178], lumberyards[1178]}), .init(2'b01), .state({trees[1127], lumberyards[1127]}));
acre acre_22_28 (.clk(clk), .en(en), .top_left({trees[1077], lumberyards[1077]}), .top({trees[1078], lumberyards[1078]}), .top_right({trees[1079], lumberyards[1079]}), .left({trees[1127], lumberyards[1127]}), .right({trees[1129], lumberyards[1129]}), .bottom_left({trees[1177], lumberyards[1177]}), .bottom({trees[1178], lumberyards[1178]}), .bottom_right({trees[1179], lumberyards[1179]}), .init(2'b10), .state({trees[1128], lumberyards[1128]}));
acre acre_22_29 (.clk(clk), .en(en), .top_left({trees[1078], lumberyards[1078]}), .top({trees[1079], lumberyards[1079]}), .top_right({trees[1080], lumberyards[1080]}), .left({trees[1128], lumberyards[1128]}), .right({trees[1130], lumberyards[1130]}), .bottom_left({trees[1178], lumberyards[1178]}), .bottom({trees[1179], lumberyards[1179]}), .bottom_right({trees[1180], lumberyards[1180]}), .init(2'b00), .state({trees[1129], lumberyards[1129]}));
acre acre_22_30 (.clk(clk), .en(en), .top_left({trees[1079], lumberyards[1079]}), .top({trees[1080], lumberyards[1080]}), .top_right({trees[1081], lumberyards[1081]}), .left({trees[1129], lumberyards[1129]}), .right({trees[1131], lumberyards[1131]}), .bottom_left({trees[1179], lumberyards[1179]}), .bottom({trees[1180], lumberyards[1180]}), .bottom_right({trees[1181], lumberyards[1181]}), .init(2'b00), .state({trees[1130], lumberyards[1130]}));
acre acre_22_31 (.clk(clk), .en(en), .top_left({trees[1080], lumberyards[1080]}), .top({trees[1081], lumberyards[1081]}), .top_right({trees[1082], lumberyards[1082]}), .left({trees[1130], lumberyards[1130]}), .right({trees[1132], lumberyards[1132]}), .bottom_left({trees[1180], lumberyards[1180]}), .bottom({trees[1181], lumberyards[1181]}), .bottom_right({trees[1182], lumberyards[1182]}), .init(2'b00), .state({trees[1131], lumberyards[1131]}));
acre acre_22_32 (.clk(clk), .en(en), .top_left({trees[1081], lumberyards[1081]}), .top({trees[1082], lumberyards[1082]}), .top_right({trees[1083], lumberyards[1083]}), .left({trees[1131], lumberyards[1131]}), .right({trees[1133], lumberyards[1133]}), .bottom_left({trees[1181], lumberyards[1181]}), .bottom({trees[1182], lumberyards[1182]}), .bottom_right({trees[1183], lumberyards[1183]}), .init(2'b01), .state({trees[1132], lumberyards[1132]}));
acre acre_22_33 (.clk(clk), .en(en), .top_left({trees[1082], lumberyards[1082]}), .top({trees[1083], lumberyards[1083]}), .top_right({trees[1084], lumberyards[1084]}), .left({trees[1132], lumberyards[1132]}), .right({trees[1134], lumberyards[1134]}), .bottom_left({trees[1182], lumberyards[1182]}), .bottom({trees[1183], lumberyards[1183]}), .bottom_right({trees[1184], lumberyards[1184]}), .init(2'b00), .state({trees[1133], lumberyards[1133]}));
acre acre_22_34 (.clk(clk), .en(en), .top_left({trees[1083], lumberyards[1083]}), .top({trees[1084], lumberyards[1084]}), .top_right({trees[1085], lumberyards[1085]}), .left({trees[1133], lumberyards[1133]}), .right({trees[1135], lumberyards[1135]}), .bottom_left({trees[1183], lumberyards[1183]}), .bottom({trees[1184], lumberyards[1184]}), .bottom_right({trees[1185], lumberyards[1185]}), .init(2'b00), .state({trees[1134], lumberyards[1134]}));
acre acre_22_35 (.clk(clk), .en(en), .top_left({trees[1084], lumberyards[1084]}), .top({trees[1085], lumberyards[1085]}), .top_right({trees[1086], lumberyards[1086]}), .left({trees[1134], lumberyards[1134]}), .right({trees[1136], lumberyards[1136]}), .bottom_left({trees[1184], lumberyards[1184]}), .bottom({trees[1185], lumberyards[1185]}), .bottom_right({trees[1186], lumberyards[1186]}), .init(2'b01), .state({trees[1135], lumberyards[1135]}));
acre acre_22_36 (.clk(clk), .en(en), .top_left({trees[1085], lumberyards[1085]}), .top({trees[1086], lumberyards[1086]}), .top_right({trees[1087], lumberyards[1087]}), .left({trees[1135], lumberyards[1135]}), .right({trees[1137], lumberyards[1137]}), .bottom_left({trees[1185], lumberyards[1185]}), .bottom({trees[1186], lumberyards[1186]}), .bottom_right({trees[1187], lumberyards[1187]}), .init(2'b01), .state({trees[1136], lumberyards[1136]}));
acre acre_22_37 (.clk(clk), .en(en), .top_left({trees[1086], lumberyards[1086]}), .top({trees[1087], lumberyards[1087]}), .top_right({trees[1088], lumberyards[1088]}), .left({trees[1136], lumberyards[1136]}), .right({trees[1138], lumberyards[1138]}), .bottom_left({trees[1186], lumberyards[1186]}), .bottom({trees[1187], lumberyards[1187]}), .bottom_right({trees[1188], lumberyards[1188]}), .init(2'b00), .state({trees[1137], lumberyards[1137]}));
acre acre_22_38 (.clk(clk), .en(en), .top_left({trees[1087], lumberyards[1087]}), .top({trees[1088], lumberyards[1088]}), .top_right({trees[1089], lumberyards[1089]}), .left({trees[1137], lumberyards[1137]}), .right({trees[1139], lumberyards[1139]}), .bottom_left({trees[1187], lumberyards[1187]}), .bottom({trees[1188], lumberyards[1188]}), .bottom_right({trees[1189], lumberyards[1189]}), .init(2'b00), .state({trees[1138], lumberyards[1138]}));
acre acre_22_39 (.clk(clk), .en(en), .top_left({trees[1088], lumberyards[1088]}), .top({trees[1089], lumberyards[1089]}), .top_right({trees[1090], lumberyards[1090]}), .left({trees[1138], lumberyards[1138]}), .right({trees[1140], lumberyards[1140]}), .bottom_left({trees[1188], lumberyards[1188]}), .bottom({trees[1189], lumberyards[1189]}), .bottom_right({trees[1190], lumberyards[1190]}), .init(2'b01), .state({trees[1139], lumberyards[1139]}));
acre acre_22_40 (.clk(clk), .en(en), .top_left({trees[1089], lumberyards[1089]}), .top({trees[1090], lumberyards[1090]}), .top_right({trees[1091], lumberyards[1091]}), .left({trees[1139], lumberyards[1139]}), .right({trees[1141], lumberyards[1141]}), .bottom_left({trees[1189], lumberyards[1189]}), .bottom({trees[1190], lumberyards[1190]}), .bottom_right({trees[1191], lumberyards[1191]}), .init(2'b00), .state({trees[1140], lumberyards[1140]}));
acre acre_22_41 (.clk(clk), .en(en), .top_left({trees[1090], lumberyards[1090]}), .top({trees[1091], lumberyards[1091]}), .top_right({trees[1092], lumberyards[1092]}), .left({trees[1140], lumberyards[1140]}), .right({trees[1142], lumberyards[1142]}), .bottom_left({trees[1190], lumberyards[1190]}), .bottom({trees[1191], lumberyards[1191]}), .bottom_right({trees[1192], lumberyards[1192]}), .init(2'b10), .state({trees[1141], lumberyards[1141]}));
acre acre_22_42 (.clk(clk), .en(en), .top_left({trees[1091], lumberyards[1091]}), .top({trees[1092], lumberyards[1092]}), .top_right({trees[1093], lumberyards[1093]}), .left({trees[1141], lumberyards[1141]}), .right({trees[1143], lumberyards[1143]}), .bottom_left({trees[1191], lumberyards[1191]}), .bottom({trees[1192], lumberyards[1192]}), .bottom_right({trees[1193], lumberyards[1193]}), .init(2'b01), .state({trees[1142], lumberyards[1142]}));
acre acre_22_43 (.clk(clk), .en(en), .top_left({trees[1092], lumberyards[1092]}), .top({trees[1093], lumberyards[1093]}), .top_right({trees[1094], lumberyards[1094]}), .left({trees[1142], lumberyards[1142]}), .right({trees[1144], lumberyards[1144]}), .bottom_left({trees[1192], lumberyards[1192]}), .bottom({trees[1193], lumberyards[1193]}), .bottom_right({trees[1194], lumberyards[1194]}), .init(2'b01), .state({trees[1143], lumberyards[1143]}));
acre acre_22_44 (.clk(clk), .en(en), .top_left({trees[1093], lumberyards[1093]}), .top({trees[1094], lumberyards[1094]}), .top_right({trees[1095], lumberyards[1095]}), .left({trees[1143], lumberyards[1143]}), .right({trees[1145], lumberyards[1145]}), .bottom_left({trees[1193], lumberyards[1193]}), .bottom({trees[1194], lumberyards[1194]}), .bottom_right({trees[1195], lumberyards[1195]}), .init(2'b00), .state({trees[1144], lumberyards[1144]}));
acre acre_22_45 (.clk(clk), .en(en), .top_left({trees[1094], lumberyards[1094]}), .top({trees[1095], lumberyards[1095]}), .top_right({trees[1096], lumberyards[1096]}), .left({trees[1144], lumberyards[1144]}), .right({trees[1146], lumberyards[1146]}), .bottom_left({trees[1194], lumberyards[1194]}), .bottom({trees[1195], lumberyards[1195]}), .bottom_right({trees[1196], lumberyards[1196]}), .init(2'b10), .state({trees[1145], lumberyards[1145]}));
acre acre_22_46 (.clk(clk), .en(en), .top_left({trees[1095], lumberyards[1095]}), .top({trees[1096], lumberyards[1096]}), .top_right({trees[1097], lumberyards[1097]}), .left({trees[1145], lumberyards[1145]}), .right({trees[1147], lumberyards[1147]}), .bottom_left({trees[1195], lumberyards[1195]}), .bottom({trees[1196], lumberyards[1196]}), .bottom_right({trees[1197], lumberyards[1197]}), .init(2'b10), .state({trees[1146], lumberyards[1146]}));
acre acre_22_47 (.clk(clk), .en(en), .top_left({trees[1096], lumberyards[1096]}), .top({trees[1097], lumberyards[1097]}), .top_right({trees[1098], lumberyards[1098]}), .left({trees[1146], lumberyards[1146]}), .right({trees[1148], lumberyards[1148]}), .bottom_left({trees[1196], lumberyards[1196]}), .bottom({trees[1197], lumberyards[1197]}), .bottom_right({trees[1198], lumberyards[1198]}), .init(2'b01), .state({trees[1147], lumberyards[1147]}));
acre acre_22_48 (.clk(clk), .en(en), .top_left({trees[1097], lumberyards[1097]}), .top({trees[1098], lumberyards[1098]}), .top_right({trees[1099], lumberyards[1099]}), .left({trees[1147], lumberyards[1147]}), .right({trees[1149], lumberyards[1149]}), .bottom_left({trees[1197], lumberyards[1197]}), .bottom({trees[1198], lumberyards[1198]}), .bottom_right({trees[1199], lumberyards[1199]}), .init(2'b01), .state({trees[1148], lumberyards[1148]}));
acre acre_22_49 (.clk(clk), .en(en), .top_left({trees[1098], lumberyards[1098]}), .top({trees[1099], lumberyards[1099]}), .top_right(2'b0), .left({trees[1148], lumberyards[1148]}), .right(2'b0), .bottom_left({trees[1198], lumberyards[1198]}), .bottom({trees[1199], lumberyards[1199]}), .bottom_right(2'b0), .init(2'b10), .state({trees[1149], lumberyards[1149]}));
acre acre_23_0 (.clk(clk), .en(en), .top_left(2'b0), .top({trees[1100], lumberyards[1100]}), .top_right({trees[1101], lumberyards[1101]}), .left(2'b0), .right({trees[1151], lumberyards[1151]}), .bottom_left(2'b0), .bottom({trees[1200], lumberyards[1200]}), .bottom_right({trees[1201], lumberyards[1201]}), .init(2'b00), .state({trees[1150], lumberyards[1150]}));
acre acre_23_1 (.clk(clk), .en(en), .top_left({trees[1100], lumberyards[1100]}), .top({trees[1101], lumberyards[1101]}), .top_right({trees[1102], lumberyards[1102]}), .left({trees[1150], lumberyards[1150]}), .right({trees[1152], lumberyards[1152]}), .bottom_left({trees[1200], lumberyards[1200]}), .bottom({trees[1201], lumberyards[1201]}), .bottom_right({trees[1202], lumberyards[1202]}), .init(2'b00), .state({trees[1151], lumberyards[1151]}));
acre acre_23_2 (.clk(clk), .en(en), .top_left({trees[1101], lumberyards[1101]}), .top({trees[1102], lumberyards[1102]}), .top_right({trees[1103], lumberyards[1103]}), .left({trees[1151], lumberyards[1151]}), .right({trees[1153], lumberyards[1153]}), .bottom_left({trees[1201], lumberyards[1201]}), .bottom({trees[1202], lumberyards[1202]}), .bottom_right({trees[1203], lumberyards[1203]}), .init(2'b10), .state({trees[1152], lumberyards[1152]}));
acre acre_23_3 (.clk(clk), .en(en), .top_left({trees[1102], lumberyards[1102]}), .top({trees[1103], lumberyards[1103]}), .top_right({trees[1104], lumberyards[1104]}), .left({trees[1152], lumberyards[1152]}), .right({trees[1154], lumberyards[1154]}), .bottom_left({trees[1202], lumberyards[1202]}), .bottom({trees[1203], lumberyards[1203]}), .bottom_right({trees[1204], lumberyards[1204]}), .init(2'b10), .state({trees[1153], lumberyards[1153]}));
acre acre_23_4 (.clk(clk), .en(en), .top_left({trees[1103], lumberyards[1103]}), .top({trees[1104], lumberyards[1104]}), .top_right({trees[1105], lumberyards[1105]}), .left({trees[1153], lumberyards[1153]}), .right({trees[1155], lumberyards[1155]}), .bottom_left({trees[1203], lumberyards[1203]}), .bottom({trees[1204], lumberyards[1204]}), .bottom_right({trees[1205], lumberyards[1205]}), .init(2'b10), .state({trees[1154], lumberyards[1154]}));
acre acre_23_5 (.clk(clk), .en(en), .top_left({trees[1104], lumberyards[1104]}), .top({trees[1105], lumberyards[1105]}), .top_right({trees[1106], lumberyards[1106]}), .left({trees[1154], lumberyards[1154]}), .right({trees[1156], lumberyards[1156]}), .bottom_left({trees[1204], lumberyards[1204]}), .bottom({trees[1205], lumberyards[1205]}), .bottom_right({trees[1206], lumberyards[1206]}), .init(2'b00), .state({trees[1155], lumberyards[1155]}));
acre acre_23_6 (.clk(clk), .en(en), .top_left({trees[1105], lumberyards[1105]}), .top({trees[1106], lumberyards[1106]}), .top_right({trees[1107], lumberyards[1107]}), .left({trees[1155], lumberyards[1155]}), .right({trees[1157], lumberyards[1157]}), .bottom_left({trees[1205], lumberyards[1205]}), .bottom({trees[1206], lumberyards[1206]}), .bottom_right({trees[1207], lumberyards[1207]}), .init(2'b00), .state({trees[1156], lumberyards[1156]}));
acre acre_23_7 (.clk(clk), .en(en), .top_left({trees[1106], lumberyards[1106]}), .top({trees[1107], lumberyards[1107]}), .top_right({trees[1108], lumberyards[1108]}), .left({trees[1156], lumberyards[1156]}), .right({trees[1158], lumberyards[1158]}), .bottom_left({trees[1206], lumberyards[1206]}), .bottom({trees[1207], lumberyards[1207]}), .bottom_right({trees[1208], lumberyards[1208]}), .init(2'b00), .state({trees[1157], lumberyards[1157]}));
acre acre_23_8 (.clk(clk), .en(en), .top_left({trees[1107], lumberyards[1107]}), .top({trees[1108], lumberyards[1108]}), .top_right({trees[1109], lumberyards[1109]}), .left({trees[1157], lumberyards[1157]}), .right({trees[1159], lumberyards[1159]}), .bottom_left({trees[1207], lumberyards[1207]}), .bottom({trees[1208], lumberyards[1208]}), .bottom_right({trees[1209], lumberyards[1209]}), .init(2'b00), .state({trees[1158], lumberyards[1158]}));
acre acre_23_9 (.clk(clk), .en(en), .top_left({trees[1108], lumberyards[1108]}), .top({trees[1109], lumberyards[1109]}), .top_right({trees[1110], lumberyards[1110]}), .left({trees[1158], lumberyards[1158]}), .right({trees[1160], lumberyards[1160]}), .bottom_left({trees[1208], lumberyards[1208]}), .bottom({trees[1209], lumberyards[1209]}), .bottom_right({trees[1210], lumberyards[1210]}), .init(2'b00), .state({trees[1159], lumberyards[1159]}));
acre acre_23_10 (.clk(clk), .en(en), .top_left({trees[1109], lumberyards[1109]}), .top({trees[1110], lumberyards[1110]}), .top_right({trees[1111], lumberyards[1111]}), .left({trees[1159], lumberyards[1159]}), .right({trees[1161], lumberyards[1161]}), .bottom_left({trees[1209], lumberyards[1209]}), .bottom({trees[1210], lumberyards[1210]}), .bottom_right({trees[1211], lumberyards[1211]}), .init(2'b00), .state({trees[1160], lumberyards[1160]}));
acre acre_23_11 (.clk(clk), .en(en), .top_left({trees[1110], lumberyards[1110]}), .top({trees[1111], lumberyards[1111]}), .top_right({trees[1112], lumberyards[1112]}), .left({trees[1160], lumberyards[1160]}), .right({trees[1162], lumberyards[1162]}), .bottom_left({trees[1210], lumberyards[1210]}), .bottom({trees[1211], lumberyards[1211]}), .bottom_right({trees[1212], lumberyards[1212]}), .init(2'b01), .state({trees[1161], lumberyards[1161]}));
acre acre_23_12 (.clk(clk), .en(en), .top_left({trees[1111], lumberyards[1111]}), .top({trees[1112], lumberyards[1112]}), .top_right({trees[1113], lumberyards[1113]}), .left({trees[1161], lumberyards[1161]}), .right({trees[1163], lumberyards[1163]}), .bottom_left({trees[1211], lumberyards[1211]}), .bottom({trees[1212], lumberyards[1212]}), .bottom_right({trees[1213], lumberyards[1213]}), .init(2'b10), .state({trees[1162], lumberyards[1162]}));
acre acre_23_13 (.clk(clk), .en(en), .top_left({trees[1112], lumberyards[1112]}), .top({trees[1113], lumberyards[1113]}), .top_right({trees[1114], lumberyards[1114]}), .left({trees[1162], lumberyards[1162]}), .right({trees[1164], lumberyards[1164]}), .bottom_left({trees[1212], lumberyards[1212]}), .bottom({trees[1213], lumberyards[1213]}), .bottom_right({trees[1214], lumberyards[1214]}), .init(2'b00), .state({trees[1163], lumberyards[1163]}));
acre acre_23_14 (.clk(clk), .en(en), .top_left({trees[1113], lumberyards[1113]}), .top({trees[1114], lumberyards[1114]}), .top_right({trees[1115], lumberyards[1115]}), .left({trees[1163], lumberyards[1163]}), .right({trees[1165], lumberyards[1165]}), .bottom_left({trees[1213], lumberyards[1213]}), .bottom({trees[1214], lumberyards[1214]}), .bottom_right({trees[1215], lumberyards[1215]}), .init(2'b00), .state({trees[1164], lumberyards[1164]}));
acre acre_23_15 (.clk(clk), .en(en), .top_left({trees[1114], lumberyards[1114]}), .top({trees[1115], lumberyards[1115]}), .top_right({trees[1116], lumberyards[1116]}), .left({trees[1164], lumberyards[1164]}), .right({trees[1166], lumberyards[1166]}), .bottom_left({trees[1214], lumberyards[1214]}), .bottom({trees[1215], lumberyards[1215]}), .bottom_right({trees[1216], lumberyards[1216]}), .init(2'b00), .state({trees[1165], lumberyards[1165]}));
acre acre_23_16 (.clk(clk), .en(en), .top_left({trees[1115], lumberyards[1115]}), .top({trees[1116], lumberyards[1116]}), .top_right({trees[1117], lumberyards[1117]}), .left({trees[1165], lumberyards[1165]}), .right({trees[1167], lumberyards[1167]}), .bottom_left({trees[1215], lumberyards[1215]}), .bottom({trees[1216], lumberyards[1216]}), .bottom_right({trees[1217], lumberyards[1217]}), .init(2'b00), .state({trees[1166], lumberyards[1166]}));
acre acre_23_17 (.clk(clk), .en(en), .top_left({trees[1116], lumberyards[1116]}), .top({trees[1117], lumberyards[1117]}), .top_right({trees[1118], lumberyards[1118]}), .left({trees[1166], lumberyards[1166]}), .right({trees[1168], lumberyards[1168]}), .bottom_left({trees[1216], lumberyards[1216]}), .bottom({trees[1217], lumberyards[1217]}), .bottom_right({trees[1218], lumberyards[1218]}), .init(2'b00), .state({trees[1167], lumberyards[1167]}));
acre acre_23_18 (.clk(clk), .en(en), .top_left({trees[1117], lumberyards[1117]}), .top({trees[1118], lumberyards[1118]}), .top_right({trees[1119], lumberyards[1119]}), .left({trees[1167], lumberyards[1167]}), .right({trees[1169], lumberyards[1169]}), .bottom_left({trees[1217], lumberyards[1217]}), .bottom({trees[1218], lumberyards[1218]}), .bottom_right({trees[1219], lumberyards[1219]}), .init(2'b00), .state({trees[1168], lumberyards[1168]}));
acre acre_23_19 (.clk(clk), .en(en), .top_left({trees[1118], lumberyards[1118]}), .top({trees[1119], lumberyards[1119]}), .top_right({trees[1120], lumberyards[1120]}), .left({trees[1168], lumberyards[1168]}), .right({trees[1170], lumberyards[1170]}), .bottom_left({trees[1218], lumberyards[1218]}), .bottom({trees[1219], lumberyards[1219]}), .bottom_right({trees[1220], lumberyards[1220]}), .init(2'b10), .state({trees[1169], lumberyards[1169]}));
acre acre_23_20 (.clk(clk), .en(en), .top_left({trees[1119], lumberyards[1119]}), .top({trees[1120], lumberyards[1120]}), .top_right({trees[1121], lumberyards[1121]}), .left({trees[1169], lumberyards[1169]}), .right({trees[1171], lumberyards[1171]}), .bottom_left({trees[1219], lumberyards[1219]}), .bottom({trees[1220], lumberyards[1220]}), .bottom_right({trees[1221], lumberyards[1221]}), .init(2'b00), .state({trees[1170], lumberyards[1170]}));
acre acre_23_21 (.clk(clk), .en(en), .top_left({trees[1120], lumberyards[1120]}), .top({trees[1121], lumberyards[1121]}), .top_right({trees[1122], lumberyards[1122]}), .left({trees[1170], lumberyards[1170]}), .right({trees[1172], lumberyards[1172]}), .bottom_left({trees[1220], lumberyards[1220]}), .bottom({trees[1221], lumberyards[1221]}), .bottom_right({trees[1222], lumberyards[1222]}), .init(2'b00), .state({trees[1171], lumberyards[1171]}));
acre acre_23_22 (.clk(clk), .en(en), .top_left({trees[1121], lumberyards[1121]}), .top({trees[1122], lumberyards[1122]}), .top_right({trees[1123], lumberyards[1123]}), .left({trees[1171], lumberyards[1171]}), .right({trees[1173], lumberyards[1173]}), .bottom_left({trees[1221], lumberyards[1221]}), .bottom({trees[1222], lumberyards[1222]}), .bottom_right({trees[1223], lumberyards[1223]}), .init(2'b10), .state({trees[1172], lumberyards[1172]}));
acre acre_23_23 (.clk(clk), .en(en), .top_left({trees[1122], lumberyards[1122]}), .top({trees[1123], lumberyards[1123]}), .top_right({trees[1124], lumberyards[1124]}), .left({trees[1172], lumberyards[1172]}), .right({trees[1174], lumberyards[1174]}), .bottom_left({trees[1222], lumberyards[1222]}), .bottom({trees[1223], lumberyards[1223]}), .bottom_right({trees[1224], lumberyards[1224]}), .init(2'b01), .state({trees[1173], lumberyards[1173]}));
acre acre_23_24 (.clk(clk), .en(en), .top_left({trees[1123], lumberyards[1123]}), .top({trees[1124], lumberyards[1124]}), .top_right({trees[1125], lumberyards[1125]}), .left({trees[1173], lumberyards[1173]}), .right({trees[1175], lumberyards[1175]}), .bottom_left({trees[1223], lumberyards[1223]}), .bottom({trees[1224], lumberyards[1224]}), .bottom_right({trees[1225], lumberyards[1225]}), .init(2'b00), .state({trees[1174], lumberyards[1174]}));
acre acre_23_25 (.clk(clk), .en(en), .top_left({trees[1124], lumberyards[1124]}), .top({trees[1125], lumberyards[1125]}), .top_right({trees[1126], lumberyards[1126]}), .left({trees[1174], lumberyards[1174]}), .right({trees[1176], lumberyards[1176]}), .bottom_left({trees[1224], lumberyards[1224]}), .bottom({trees[1225], lumberyards[1225]}), .bottom_right({trees[1226], lumberyards[1226]}), .init(2'b10), .state({trees[1175], lumberyards[1175]}));
acre acre_23_26 (.clk(clk), .en(en), .top_left({trees[1125], lumberyards[1125]}), .top({trees[1126], lumberyards[1126]}), .top_right({trees[1127], lumberyards[1127]}), .left({trees[1175], lumberyards[1175]}), .right({trees[1177], lumberyards[1177]}), .bottom_left({trees[1225], lumberyards[1225]}), .bottom({trees[1226], lumberyards[1226]}), .bottom_right({trees[1227], lumberyards[1227]}), .init(2'b10), .state({trees[1176], lumberyards[1176]}));
acre acre_23_27 (.clk(clk), .en(en), .top_left({trees[1126], lumberyards[1126]}), .top({trees[1127], lumberyards[1127]}), .top_right({trees[1128], lumberyards[1128]}), .left({trees[1176], lumberyards[1176]}), .right({trees[1178], lumberyards[1178]}), .bottom_left({trees[1226], lumberyards[1226]}), .bottom({trees[1227], lumberyards[1227]}), .bottom_right({trees[1228], lumberyards[1228]}), .init(2'b00), .state({trees[1177], lumberyards[1177]}));
acre acre_23_28 (.clk(clk), .en(en), .top_left({trees[1127], lumberyards[1127]}), .top({trees[1128], lumberyards[1128]}), .top_right({trees[1129], lumberyards[1129]}), .left({trees[1177], lumberyards[1177]}), .right({trees[1179], lumberyards[1179]}), .bottom_left({trees[1227], lumberyards[1227]}), .bottom({trees[1228], lumberyards[1228]}), .bottom_right({trees[1229], lumberyards[1229]}), .init(2'b10), .state({trees[1178], lumberyards[1178]}));
acre acre_23_29 (.clk(clk), .en(en), .top_left({trees[1128], lumberyards[1128]}), .top({trees[1129], lumberyards[1129]}), .top_right({trees[1130], lumberyards[1130]}), .left({trees[1178], lumberyards[1178]}), .right({trees[1180], lumberyards[1180]}), .bottom_left({trees[1228], lumberyards[1228]}), .bottom({trees[1229], lumberyards[1229]}), .bottom_right({trees[1230], lumberyards[1230]}), .init(2'b01), .state({trees[1179], lumberyards[1179]}));
acre acre_23_30 (.clk(clk), .en(en), .top_left({trees[1129], lumberyards[1129]}), .top({trees[1130], lumberyards[1130]}), .top_right({trees[1131], lumberyards[1131]}), .left({trees[1179], lumberyards[1179]}), .right({trees[1181], lumberyards[1181]}), .bottom_left({trees[1229], lumberyards[1229]}), .bottom({trees[1230], lumberyards[1230]}), .bottom_right({trees[1231], lumberyards[1231]}), .init(2'b00), .state({trees[1180], lumberyards[1180]}));
acre acre_23_31 (.clk(clk), .en(en), .top_left({trees[1130], lumberyards[1130]}), .top({trees[1131], lumberyards[1131]}), .top_right({trees[1132], lumberyards[1132]}), .left({trees[1180], lumberyards[1180]}), .right({trees[1182], lumberyards[1182]}), .bottom_left({trees[1230], lumberyards[1230]}), .bottom({trees[1231], lumberyards[1231]}), .bottom_right({trees[1232], lumberyards[1232]}), .init(2'b10), .state({trees[1181], lumberyards[1181]}));
acre acre_23_32 (.clk(clk), .en(en), .top_left({trees[1131], lumberyards[1131]}), .top({trees[1132], lumberyards[1132]}), .top_right({trees[1133], lumberyards[1133]}), .left({trees[1181], lumberyards[1181]}), .right({trees[1183], lumberyards[1183]}), .bottom_left({trees[1231], lumberyards[1231]}), .bottom({trees[1232], lumberyards[1232]}), .bottom_right({trees[1233], lumberyards[1233]}), .init(2'b01), .state({trees[1182], lumberyards[1182]}));
acre acre_23_33 (.clk(clk), .en(en), .top_left({trees[1132], lumberyards[1132]}), .top({trees[1133], lumberyards[1133]}), .top_right({trees[1134], lumberyards[1134]}), .left({trees[1182], lumberyards[1182]}), .right({trees[1184], lumberyards[1184]}), .bottom_left({trees[1232], lumberyards[1232]}), .bottom({trees[1233], lumberyards[1233]}), .bottom_right({trees[1234], lumberyards[1234]}), .init(2'b00), .state({trees[1183], lumberyards[1183]}));
acre acre_23_34 (.clk(clk), .en(en), .top_left({trees[1133], lumberyards[1133]}), .top({trees[1134], lumberyards[1134]}), .top_right({trees[1135], lumberyards[1135]}), .left({trees[1183], lumberyards[1183]}), .right({trees[1185], lumberyards[1185]}), .bottom_left({trees[1233], lumberyards[1233]}), .bottom({trees[1234], lumberyards[1234]}), .bottom_right({trees[1235], lumberyards[1235]}), .init(2'b00), .state({trees[1184], lumberyards[1184]}));
acre acre_23_35 (.clk(clk), .en(en), .top_left({trees[1134], lumberyards[1134]}), .top({trees[1135], lumberyards[1135]}), .top_right({trees[1136], lumberyards[1136]}), .left({trees[1184], lumberyards[1184]}), .right({trees[1186], lumberyards[1186]}), .bottom_left({trees[1234], lumberyards[1234]}), .bottom({trees[1235], lumberyards[1235]}), .bottom_right({trees[1236], lumberyards[1236]}), .init(2'b01), .state({trees[1185], lumberyards[1185]}));
acre acre_23_36 (.clk(clk), .en(en), .top_left({trees[1135], lumberyards[1135]}), .top({trees[1136], lumberyards[1136]}), .top_right({trees[1137], lumberyards[1137]}), .left({trees[1185], lumberyards[1185]}), .right({trees[1187], lumberyards[1187]}), .bottom_left({trees[1235], lumberyards[1235]}), .bottom({trees[1236], lumberyards[1236]}), .bottom_right({trees[1237], lumberyards[1237]}), .init(2'b00), .state({trees[1186], lumberyards[1186]}));
acre acre_23_37 (.clk(clk), .en(en), .top_left({trees[1136], lumberyards[1136]}), .top({trees[1137], lumberyards[1137]}), .top_right({trees[1138], lumberyards[1138]}), .left({trees[1186], lumberyards[1186]}), .right({trees[1188], lumberyards[1188]}), .bottom_left({trees[1236], lumberyards[1236]}), .bottom({trees[1237], lumberyards[1237]}), .bottom_right({trees[1238], lumberyards[1238]}), .init(2'b00), .state({trees[1187], lumberyards[1187]}));
acre acre_23_38 (.clk(clk), .en(en), .top_left({trees[1137], lumberyards[1137]}), .top({trees[1138], lumberyards[1138]}), .top_right({trees[1139], lumberyards[1139]}), .left({trees[1187], lumberyards[1187]}), .right({trees[1189], lumberyards[1189]}), .bottom_left({trees[1237], lumberyards[1237]}), .bottom({trees[1238], lumberyards[1238]}), .bottom_right({trees[1239], lumberyards[1239]}), .init(2'b00), .state({trees[1188], lumberyards[1188]}));
acre acre_23_39 (.clk(clk), .en(en), .top_left({trees[1138], lumberyards[1138]}), .top({trees[1139], lumberyards[1139]}), .top_right({trees[1140], lumberyards[1140]}), .left({trees[1188], lumberyards[1188]}), .right({trees[1190], lumberyards[1190]}), .bottom_left({trees[1238], lumberyards[1238]}), .bottom({trees[1239], lumberyards[1239]}), .bottom_right({trees[1240], lumberyards[1240]}), .init(2'b01), .state({trees[1189], lumberyards[1189]}));
acre acre_23_40 (.clk(clk), .en(en), .top_left({trees[1139], lumberyards[1139]}), .top({trees[1140], lumberyards[1140]}), .top_right({trees[1141], lumberyards[1141]}), .left({trees[1189], lumberyards[1189]}), .right({trees[1191], lumberyards[1191]}), .bottom_left({trees[1239], lumberyards[1239]}), .bottom({trees[1240], lumberyards[1240]}), .bottom_right({trees[1241], lumberyards[1241]}), .init(2'b00), .state({trees[1190], lumberyards[1190]}));
acre acre_23_41 (.clk(clk), .en(en), .top_left({trees[1140], lumberyards[1140]}), .top({trees[1141], lumberyards[1141]}), .top_right({trees[1142], lumberyards[1142]}), .left({trees[1190], lumberyards[1190]}), .right({trees[1192], lumberyards[1192]}), .bottom_left({trees[1240], lumberyards[1240]}), .bottom({trees[1241], lumberyards[1241]}), .bottom_right({trees[1242], lumberyards[1242]}), .init(2'b10), .state({trees[1191], lumberyards[1191]}));
acre acre_23_42 (.clk(clk), .en(en), .top_left({trees[1141], lumberyards[1141]}), .top({trees[1142], lumberyards[1142]}), .top_right({trees[1143], lumberyards[1143]}), .left({trees[1191], lumberyards[1191]}), .right({trees[1193], lumberyards[1193]}), .bottom_left({trees[1241], lumberyards[1241]}), .bottom({trees[1242], lumberyards[1242]}), .bottom_right({trees[1243], lumberyards[1243]}), .init(2'b00), .state({trees[1192], lumberyards[1192]}));
acre acre_23_43 (.clk(clk), .en(en), .top_left({trees[1142], lumberyards[1142]}), .top({trees[1143], lumberyards[1143]}), .top_right({trees[1144], lumberyards[1144]}), .left({trees[1192], lumberyards[1192]}), .right({trees[1194], lumberyards[1194]}), .bottom_left({trees[1242], lumberyards[1242]}), .bottom({trees[1243], lumberyards[1243]}), .bottom_right({trees[1244], lumberyards[1244]}), .init(2'b10), .state({trees[1193], lumberyards[1193]}));
acre acre_23_44 (.clk(clk), .en(en), .top_left({trees[1143], lumberyards[1143]}), .top({trees[1144], lumberyards[1144]}), .top_right({trees[1145], lumberyards[1145]}), .left({trees[1193], lumberyards[1193]}), .right({trees[1195], lumberyards[1195]}), .bottom_left({trees[1243], lumberyards[1243]}), .bottom({trees[1244], lumberyards[1244]}), .bottom_right({trees[1245], lumberyards[1245]}), .init(2'b00), .state({trees[1194], lumberyards[1194]}));
acre acre_23_45 (.clk(clk), .en(en), .top_left({trees[1144], lumberyards[1144]}), .top({trees[1145], lumberyards[1145]}), .top_right({trees[1146], lumberyards[1146]}), .left({trees[1194], lumberyards[1194]}), .right({trees[1196], lumberyards[1196]}), .bottom_left({trees[1244], lumberyards[1244]}), .bottom({trees[1245], lumberyards[1245]}), .bottom_right({trees[1246], lumberyards[1246]}), .init(2'b00), .state({trees[1195], lumberyards[1195]}));
acre acre_23_46 (.clk(clk), .en(en), .top_left({trees[1145], lumberyards[1145]}), .top({trees[1146], lumberyards[1146]}), .top_right({trees[1147], lumberyards[1147]}), .left({trees[1195], lumberyards[1195]}), .right({trees[1197], lumberyards[1197]}), .bottom_left({trees[1245], lumberyards[1245]}), .bottom({trees[1246], lumberyards[1246]}), .bottom_right({trees[1247], lumberyards[1247]}), .init(2'b00), .state({trees[1196], lumberyards[1196]}));
acre acre_23_47 (.clk(clk), .en(en), .top_left({trees[1146], lumberyards[1146]}), .top({trees[1147], lumberyards[1147]}), .top_right({trees[1148], lumberyards[1148]}), .left({trees[1196], lumberyards[1196]}), .right({trees[1198], lumberyards[1198]}), .bottom_left({trees[1246], lumberyards[1246]}), .bottom({trees[1247], lumberyards[1247]}), .bottom_right({trees[1248], lumberyards[1248]}), .init(2'b00), .state({trees[1197], lumberyards[1197]}));
acre acre_23_48 (.clk(clk), .en(en), .top_left({trees[1147], lumberyards[1147]}), .top({trees[1148], lumberyards[1148]}), .top_right({trees[1149], lumberyards[1149]}), .left({trees[1197], lumberyards[1197]}), .right({trees[1199], lumberyards[1199]}), .bottom_left({trees[1247], lumberyards[1247]}), .bottom({trees[1248], lumberyards[1248]}), .bottom_right({trees[1249], lumberyards[1249]}), .init(2'b00), .state({trees[1198], lumberyards[1198]}));
acre acre_23_49 (.clk(clk), .en(en), .top_left({trees[1148], lumberyards[1148]}), .top({trees[1149], lumberyards[1149]}), .top_right(2'b0), .left({trees[1198], lumberyards[1198]}), .right(2'b0), .bottom_left({trees[1248], lumberyards[1248]}), .bottom({trees[1249], lumberyards[1249]}), .bottom_right(2'b0), .init(2'b00), .state({trees[1199], lumberyards[1199]}));
acre acre_24_0 (.clk(clk), .en(en), .top_left(2'b0), .top({trees[1150], lumberyards[1150]}), .top_right({trees[1151], lumberyards[1151]}), .left(2'b0), .right({trees[1201], lumberyards[1201]}), .bottom_left(2'b0), .bottom({trees[1250], lumberyards[1250]}), .bottom_right({trees[1251], lumberyards[1251]}), .init(2'b00), .state({trees[1200], lumberyards[1200]}));
acre acre_24_1 (.clk(clk), .en(en), .top_left({trees[1150], lumberyards[1150]}), .top({trees[1151], lumberyards[1151]}), .top_right({trees[1152], lumberyards[1152]}), .left({trees[1200], lumberyards[1200]}), .right({trees[1202], lumberyards[1202]}), .bottom_left({trees[1250], lumberyards[1250]}), .bottom({trees[1251], lumberyards[1251]}), .bottom_right({trees[1252], lumberyards[1252]}), .init(2'b10), .state({trees[1201], lumberyards[1201]}));
acre acre_24_2 (.clk(clk), .en(en), .top_left({trees[1151], lumberyards[1151]}), .top({trees[1152], lumberyards[1152]}), .top_right({trees[1153], lumberyards[1153]}), .left({trees[1201], lumberyards[1201]}), .right({trees[1203], lumberyards[1203]}), .bottom_left({trees[1251], lumberyards[1251]}), .bottom({trees[1252], lumberyards[1252]}), .bottom_right({trees[1253], lumberyards[1253]}), .init(2'b00), .state({trees[1202], lumberyards[1202]}));
acre acre_24_3 (.clk(clk), .en(en), .top_left({trees[1152], lumberyards[1152]}), .top({trees[1153], lumberyards[1153]}), .top_right({trees[1154], lumberyards[1154]}), .left({trees[1202], lumberyards[1202]}), .right({trees[1204], lumberyards[1204]}), .bottom_left({trees[1252], lumberyards[1252]}), .bottom({trees[1253], lumberyards[1253]}), .bottom_right({trees[1254], lumberyards[1254]}), .init(2'b10), .state({trees[1203], lumberyards[1203]}));
acre acre_24_4 (.clk(clk), .en(en), .top_left({trees[1153], lumberyards[1153]}), .top({trees[1154], lumberyards[1154]}), .top_right({trees[1155], lumberyards[1155]}), .left({trees[1203], lumberyards[1203]}), .right({trees[1205], lumberyards[1205]}), .bottom_left({trees[1253], lumberyards[1253]}), .bottom({trees[1254], lumberyards[1254]}), .bottom_right({trees[1255], lumberyards[1255]}), .init(2'b00), .state({trees[1204], lumberyards[1204]}));
acre acre_24_5 (.clk(clk), .en(en), .top_left({trees[1154], lumberyards[1154]}), .top({trees[1155], lumberyards[1155]}), .top_right({trees[1156], lumberyards[1156]}), .left({trees[1204], lumberyards[1204]}), .right({trees[1206], lumberyards[1206]}), .bottom_left({trees[1254], lumberyards[1254]}), .bottom({trees[1255], lumberyards[1255]}), .bottom_right({trees[1256], lumberyards[1256]}), .init(2'b00), .state({trees[1205], lumberyards[1205]}));
acre acre_24_6 (.clk(clk), .en(en), .top_left({trees[1155], lumberyards[1155]}), .top({trees[1156], lumberyards[1156]}), .top_right({trees[1157], lumberyards[1157]}), .left({trees[1205], lumberyards[1205]}), .right({trees[1207], lumberyards[1207]}), .bottom_left({trees[1255], lumberyards[1255]}), .bottom({trees[1256], lumberyards[1256]}), .bottom_right({trees[1257], lumberyards[1257]}), .init(2'b01), .state({trees[1206], lumberyards[1206]}));
acre acre_24_7 (.clk(clk), .en(en), .top_left({trees[1156], lumberyards[1156]}), .top({trees[1157], lumberyards[1157]}), .top_right({trees[1158], lumberyards[1158]}), .left({trees[1206], lumberyards[1206]}), .right({trees[1208], lumberyards[1208]}), .bottom_left({trees[1256], lumberyards[1256]}), .bottom({trees[1257], lumberyards[1257]}), .bottom_right({trees[1258], lumberyards[1258]}), .init(2'b00), .state({trees[1207], lumberyards[1207]}));
acre acre_24_8 (.clk(clk), .en(en), .top_left({trees[1157], lumberyards[1157]}), .top({trees[1158], lumberyards[1158]}), .top_right({trees[1159], lumberyards[1159]}), .left({trees[1207], lumberyards[1207]}), .right({trees[1209], lumberyards[1209]}), .bottom_left({trees[1257], lumberyards[1257]}), .bottom({trees[1258], lumberyards[1258]}), .bottom_right({trees[1259], lumberyards[1259]}), .init(2'b01), .state({trees[1208], lumberyards[1208]}));
acre acre_24_9 (.clk(clk), .en(en), .top_left({trees[1158], lumberyards[1158]}), .top({trees[1159], lumberyards[1159]}), .top_right({trees[1160], lumberyards[1160]}), .left({trees[1208], lumberyards[1208]}), .right({trees[1210], lumberyards[1210]}), .bottom_left({trees[1258], lumberyards[1258]}), .bottom({trees[1259], lumberyards[1259]}), .bottom_right({trees[1260], lumberyards[1260]}), .init(2'b00), .state({trees[1209], lumberyards[1209]}));
acre acre_24_10 (.clk(clk), .en(en), .top_left({trees[1159], lumberyards[1159]}), .top({trees[1160], lumberyards[1160]}), .top_right({trees[1161], lumberyards[1161]}), .left({trees[1209], lumberyards[1209]}), .right({trees[1211], lumberyards[1211]}), .bottom_left({trees[1259], lumberyards[1259]}), .bottom({trees[1260], lumberyards[1260]}), .bottom_right({trees[1261], lumberyards[1261]}), .init(2'b01), .state({trees[1210], lumberyards[1210]}));
acre acre_24_11 (.clk(clk), .en(en), .top_left({trees[1160], lumberyards[1160]}), .top({trees[1161], lumberyards[1161]}), .top_right({trees[1162], lumberyards[1162]}), .left({trees[1210], lumberyards[1210]}), .right({trees[1212], lumberyards[1212]}), .bottom_left({trees[1260], lumberyards[1260]}), .bottom({trees[1261], lumberyards[1261]}), .bottom_right({trees[1262], lumberyards[1262]}), .init(2'b01), .state({trees[1211], lumberyards[1211]}));
acre acre_24_12 (.clk(clk), .en(en), .top_left({trees[1161], lumberyards[1161]}), .top({trees[1162], lumberyards[1162]}), .top_right({trees[1163], lumberyards[1163]}), .left({trees[1211], lumberyards[1211]}), .right({trees[1213], lumberyards[1213]}), .bottom_left({trees[1261], lumberyards[1261]}), .bottom({trees[1262], lumberyards[1262]}), .bottom_right({trees[1263], lumberyards[1263]}), .init(2'b01), .state({trees[1212], lumberyards[1212]}));
acre acre_24_13 (.clk(clk), .en(en), .top_left({trees[1162], lumberyards[1162]}), .top({trees[1163], lumberyards[1163]}), .top_right({trees[1164], lumberyards[1164]}), .left({trees[1212], lumberyards[1212]}), .right({trees[1214], lumberyards[1214]}), .bottom_left({trees[1262], lumberyards[1262]}), .bottom({trees[1263], lumberyards[1263]}), .bottom_right({trees[1264], lumberyards[1264]}), .init(2'b00), .state({trees[1213], lumberyards[1213]}));
acre acre_24_14 (.clk(clk), .en(en), .top_left({trees[1163], lumberyards[1163]}), .top({trees[1164], lumberyards[1164]}), .top_right({trees[1165], lumberyards[1165]}), .left({trees[1213], lumberyards[1213]}), .right({trees[1215], lumberyards[1215]}), .bottom_left({trees[1263], lumberyards[1263]}), .bottom({trees[1264], lumberyards[1264]}), .bottom_right({trees[1265], lumberyards[1265]}), .init(2'b00), .state({trees[1214], lumberyards[1214]}));
acre acre_24_15 (.clk(clk), .en(en), .top_left({trees[1164], lumberyards[1164]}), .top({trees[1165], lumberyards[1165]}), .top_right({trees[1166], lumberyards[1166]}), .left({trees[1214], lumberyards[1214]}), .right({trees[1216], lumberyards[1216]}), .bottom_left({trees[1264], lumberyards[1264]}), .bottom({trees[1265], lumberyards[1265]}), .bottom_right({trees[1266], lumberyards[1266]}), .init(2'b01), .state({trees[1215], lumberyards[1215]}));
acre acre_24_16 (.clk(clk), .en(en), .top_left({trees[1165], lumberyards[1165]}), .top({trees[1166], lumberyards[1166]}), .top_right({trees[1167], lumberyards[1167]}), .left({trees[1215], lumberyards[1215]}), .right({trees[1217], lumberyards[1217]}), .bottom_left({trees[1265], lumberyards[1265]}), .bottom({trees[1266], lumberyards[1266]}), .bottom_right({trees[1267], lumberyards[1267]}), .init(2'b00), .state({trees[1216], lumberyards[1216]}));
acre acre_24_17 (.clk(clk), .en(en), .top_left({trees[1166], lumberyards[1166]}), .top({trees[1167], lumberyards[1167]}), .top_right({trees[1168], lumberyards[1168]}), .left({trees[1216], lumberyards[1216]}), .right({trees[1218], lumberyards[1218]}), .bottom_left({trees[1266], lumberyards[1266]}), .bottom({trees[1267], lumberyards[1267]}), .bottom_right({trees[1268], lumberyards[1268]}), .init(2'b00), .state({trees[1217], lumberyards[1217]}));
acre acre_24_18 (.clk(clk), .en(en), .top_left({trees[1167], lumberyards[1167]}), .top({trees[1168], lumberyards[1168]}), .top_right({trees[1169], lumberyards[1169]}), .left({trees[1217], lumberyards[1217]}), .right({trees[1219], lumberyards[1219]}), .bottom_left({trees[1267], lumberyards[1267]}), .bottom({trees[1268], lumberyards[1268]}), .bottom_right({trees[1269], lumberyards[1269]}), .init(2'b01), .state({trees[1218], lumberyards[1218]}));
acre acre_24_19 (.clk(clk), .en(en), .top_left({trees[1168], lumberyards[1168]}), .top({trees[1169], lumberyards[1169]}), .top_right({trees[1170], lumberyards[1170]}), .left({trees[1218], lumberyards[1218]}), .right({trees[1220], lumberyards[1220]}), .bottom_left({trees[1268], lumberyards[1268]}), .bottom({trees[1269], lumberyards[1269]}), .bottom_right({trees[1270], lumberyards[1270]}), .init(2'b00), .state({trees[1219], lumberyards[1219]}));
acre acre_24_20 (.clk(clk), .en(en), .top_left({trees[1169], lumberyards[1169]}), .top({trees[1170], lumberyards[1170]}), .top_right({trees[1171], lumberyards[1171]}), .left({trees[1219], lumberyards[1219]}), .right({trees[1221], lumberyards[1221]}), .bottom_left({trees[1269], lumberyards[1269]}), .bottom({trees[1270], lumberyards[1270]}), .bottom_right({trees[1271], lumberyards[1271]}), .init(2'b00), .state({trees[1220], lumberyards[1220]}));
acre acre_24_21 (.clk(clk), .en(en), .top_left({trees[1170], lumberyards[1170]}), .top({trees[1171], lumberyards[1171]}), .top_right({trees[1172], lumberyards[1172]}), .left({trees[1220], lumberyards[1220]}), .right({trees[1222], lumberyards[1222]}), .bottom_left({trees[1270], lumberyards[1270]}), .bottom({trees[1271], lumberyards[1271]}), .bottom_right({trees[1272], lumberyards[1272]}), .init(2'b10), .state({trees[1221], lumberyards[1221]}));
acre acre_24_22 (.clk(clk), .en(en), .top_left({trees[1171], lumberyards[1171]}), .top({trees[1172], lumberyards[1172]}), .top_right({trees[1173], lumberyards[1173]}), .left({trees[1221], lumberyards[1221]}), .right({trees[1223], lumberyards[1223]}), .bottom_left({trees[1271], lumberyards[1271]}), .bottom({trees[1272], lumberyards[1272]}), .bottom_right({trees[1273], lumberyards[1273]}), .init(2'b01), .state({trees[1222], lumberyards[1222]}));
acre acre_24_23 (.clk(clk), .en(en), .top_left({trees[1172], lumberyards[1172]}), .top({trees[1173], lumberyards[1173]}), .top_right({trees[1174], lumberyards[1174]}), .left({trees[1222], lumberyards[1222]}), .right({trees[1224], lumberyards[1224]}), .bottom_left({trees[1272], lumberyards[1272]}), .bottom({trees[1273], lumberyards[1273]}), .bottom_right({trees[1274], lumberyards[1274]}), .init(2'b00), .state({trees[1223], lumberyards[1223]}));
acre acre_24_24 (.clk(clk), .en(en), .top_left({trees[1173], lumberyards[1173]}), .top({trees[1174], lumberyards[1174]}), .top_right({trees[1175], lumberyards[1175]}), .left({trees[1223], lumberyards[1223]}), .right({trees[1225], lumberyards[1225]}), .bottom_left({trees[1273], lumberyards[1273]}), .bottom({trees[1274], lumberyards[1274]}), .bottom_right({trees[1275], lumberyards[1275]}), .init(2'b00), .state({trees[1224], lumberyards[1224]}));
acre acre_24_25 (.clk(clk), .en(en), .top_left({trees[1174], lumberyards[1174]}), .top({trees[1175], lumberyards[1175]}), .top_right({trees[1176], lumberyards[1176]}), .left({trees[1224], lumberyards[1224]}), .right({trees[1226], lumberyards[1226]}), .bottom_left({trees[1274], lumberyards[1274]}), .bottom({trees[1275], lumberyards[1275]}), .bottom_right({trees[1276], lumberyards[1276]}), .init(2'b01), .state({trees[1225], lumberyards[1225]}));
acre acre_24_26 (.clk(clk), .en(en), .top_left({trees[1175], lumberyards[1175]}), .top({trees[1176], lumberyards[1176]}), .top_right({trees[1177], lumberyards[1177]}), .left({trees[1225], lumberyards[1225]}), .right({trees[1227], lumberyards[1227]}), .bottom_left({trees[1275], lumberyards[1275]}), .bottom({trees[1276], lumberyards[1276]}), .bottom_right({trees[1277], lumberyards[1277]}), .init(2'b00), .state({trees[1226], lumberyards[1226]}));
acre acre_24_27 (.clk(clk), .en(en), .top_left({trees[1176], lumberyards[1176]}), .top({trees[1177], lumberyards[1177]}), .top_right({trees[1178], lumberyards[1178]}), .left({trees[1226], lumberyards[1226]}), .right({trees[1228], lumberyards[1228]}), .bottom_left({trees[1276], lumberyards[1276]}), .bottom({trees[1277], lumberyards[1277]}), .bottom_right({trees[1278], lumberyards[1278]}), .init(2'b00), .state({trees[1227], lumberyards[1227]}));
acre acre_24_28 (.clk(clk), .en(en), .top_left({trees[1177], lumberyards[1177]}), .top({trees[1178], lumberyards[1178]}), .top_right({trees[1179], lumberyards[1179]}), .left({trees[1227], lumberyards[1227]}), .right({trees[1229], lumberyards[1229]}), .bottom_left({trees[1277], lumberyards[1277]}), .bottom({trees[1278], lumberyards[1278]}), .bottom_right({trees[1279], lumberyards[1279]}), .init(2'b10), .state({trees[1228], lumberyards[1228]}));
acre acre_24_29 (.clk(clk), .en(en), .top_left({trees[1178], lumberyards[1178]}), .top({trees[1179], lumberyards[1179]}), .top_right({trees[1180], lumberyards[1180]}), .left({trees[1228], lumberyards[1228]}), .right({trees[1230], lumberyards[1230]}), .bottom_left({trees[1278], lumberyards[1278]}), .bottom({trees[1279], lumberyards[1279]}), .bottom_right({trees[1280], lumberyards[1280]}), .init(2'b00), .state({trees[1229], lumberyards[1229]}));
acre acre_24_30 (.clk(clk), .en(en), .top_left({trees[1179], lumberyards[1179]}), .top({trees[1180], lumberyards[1180]}), .top_right({trees[1181], lumberyards[1181]}), .left({trees[1229], lumberyards[1229]}), .right({trees[1231], lumberyards[1231]}), .bottom_left({trees[1279], lumberyards[1279]}), .bottom({trees[1280], lumberyards[1280]}), .bottom_right({trees[1281], lumberyards[1281]}), .init(2'b00), .state({trees[1230], lumberyards[1230]}));
acre acre_24_31 (.clk(clk), .en(en), .top_left({trees[1180], lumberyards[1180]}), .top({trees[1181], lumberyards[1181]}), .top_right({trees[1182], lumberyards[1182]}), .left({trees[1230], lumberyards[1230]}), .right({trees[1232], lumberyards[1232]}), .bottom_left({trees[1280], lumberyards[1280]}), .bottom({trees[1281], lumberyards[1281]}), .bottom_right({trees[1282], lumberyards[1282]}), .init(2'b00), .state({trees[1231], lumberyards[1231]}));
acre acre_24_32 (.clk(clk), .en(en), .top_left({trees[1181], lumberyards[1181]}), .top({trees[1182], lumberyards[1182]}), .top_right({trees[1183], lumberyards[1183]}), .left({trees[1231], lumberyards[1231]}), .right({trees[1233], lumberyards[1233]}), .bottom_left({trees[1281], lumberyards[1281]}), .bottom({trees[1282], lumberyards[1282]}), .bottom_right({trees[1283], lumberyards[1283]}), .init(2'b10), .state({trees[1232], lumberyards[1232]}));
acre acre_24_33 (.clk(clk), .en(en), .top_left({trees[1182], lumberyards[1182]}), .top({trees[1183], lumberyards[1183]}), .top_right({trees[1184], lumberyards[1184]}), .left({trees[1232], lumberyards[1232]}), .right({trees[1234], lumberyards[1234]}), .bottom_left({trees[1282], lumberyards[1282]}), .bottom({trees[1283], lumberyards[1283]}), .bottom_right({trees[1284], lumberyards[1284]}), .init(2'b00), .state({trees[1233], lumberyards[1233]}));
acre acre_24_34 (.clk(clk), .en(en), .top_left({trees[1183], lumberyards[1183]}), .top({trees[1184], lumberyards[1184]}), .top_right({trees[1185], lumberyards[1185]}), .left({trees[1233], lumberyards[1233]}), .right({trees[1235], lumberyards[1235]}), .bottom_left({trees[1283], lumberyards[1283]}), .bottom({trees[1284], lumberyards[1284]}), .bottom_right({trees[1285], lumberyards[1285]}), .init(2'b00), .state({trees[1234], lumberyards[1234]}));
acre acre_24_35 (.clk(clk), .en(en), .top_left({trees[1184], lumberyards[1184]}), .top({trees[1185], lumberyards[1185]}), .top_right({trees[1186], lumberyards[1186]}), .left({trees[1234], lumberyards[1234]}), .right({trees[1236], lumberyards[1236]}), .bottom_left({trees[1284], lumberyards[1284]}), .bottom({trees[1285], lumberyards[1285]}), .bottom_right({trees[1286], lumberyards[1286]}), .init(2'b01), .state({trees[1235], lumberyards[1235]}));
acre acre_24_36 (.clk(clk), .en(en), .top_left({trees[1185], lumberyards[1185]}), .top({trees[1186], lumberyards[1186]}), .top_right({trees[1187], lumberyards[1187]}), .left({trees[1235], lumberyards[1235]}), .right({trees[1237], lumberyards[1237]}), .bottom_left({trees[1285], lumberyards[1285]}), .bottom({trees[1286], lumberyards[1286]}), .bottom_right({trees[1287], lumberyards[1287]}), .init(2'b10), .state({trees[1236], lumberyards[1236]}));
acre acre_24_37 (.clk(clk), .en(en), .top_left({trees[1186], lumberyards[1186]}), .top({trees[1187], lumberyards[1187]}), .top_right({trees[1188], lumberyards[1188]}), .left({trees[1236], lumberyards[1236]}), .right({trees[1238], lumberyards[1238]}), .bottom_left({trees[1286], lumberyards[1286]}), .bottom({trees[1287], lumberyards[1287]}), .bottom_right({trees[1288], lumberyards[1288]}), .init(2'b00), .state({trees[1237], lumberyards[1237]}));
acre acre_24_38 (.clk(clk), .en(en), .top_left({trees[1187], lumberyards[1187]}), .top({trees[1188], lumberyards[1188]}), .top_right({trees[1189], lumberyards[1189]}), .left({trees[1237], lumberyards[1237]}), .right({trees[1239], lumberyards[1239]}), .bottom_left({trees[1287], lumberyards[1287]}), .bottom({trees[1288], lumberyards[1288]}), .bottom_right({trees[1289], lumberyards[1289]}), .init(2'b00), .state({trees[1238], lumberyards[1238]}));
acre acre_24_39 (.clk(clk), .en(en), .top_left({trees[1188], lumberyards[1188]}), .top({trees[1189], lumberyards[1189]}), .top_right({trees[1190], lumberyards[1190]}), .left({trees[1238], lumberyards[1238]}), .right({trees[1240], lumberyards[1240]}), .bottom_left({trees[1288], lumberyards[1288]}), .bottom({trees[1289], lumberyards[1289]}), .bottom_right({trees[1290], lumberyards[1290]}), .init(2'b00), .state({trees[1239], lumberyards[1239]}));
acre acre_24_40 (.clk(clk), .en(en), .top_left({trees[1189], lumberyards[1189]}), .top({trees[1190], lumberyards[1190]}), .top_right({trees[1191], lumberyards[1191]}), .left({trees[1239], lumberyards[1239]}), .right({trees[1241], lumberyards[1241]}), .bottom_left({trees[1289], lumberyards[1289]}), .bottom({trees[1290], lumberyards[1290]}), .bottom_right({trees[1291], lumberyards[1291]}), .init(2'b01), .state({trees[1240], lumberyards[1240]}));
acre acre_24_41 (.clk(clk), .en(en), .top_left({trees[1190], lumberyards[1190]}), .top({trees[1191], lumberyards[1191]}), .top_right({trees[1192], lumberyards[1192]}), .left({trees[1240], lumberyards[1240]}), .right({trees[1242], lumberyards[1242]}), .bottom_left({trees[1290], lumberyards[1290]}), .bottom({trees[1291], lumberyards[1291]}), .bottom_right({trees[1292], lumberyards[1292]}), .init(2'b00), .state({trees[1241], lumberyards[1241]}));
acre acre_24_42 (.clk(clk), .en(en), .top_left({trees[1191], lumberyards[1191]}), .top({trees[1192], lumberyards[1192]}), .top_right({trees[1193], lumberyards[1193]}), .left({trees[1241], lumberyards[1241]}), .right({trees[1243], lumberyards[1243]}), .bottom_left({trees[1291], lumberyards[1291]}), .bottom({trees[1292], lumberyards[1292]}), .bottom_right({trees[1293], lumberyards[1293]}), .init(2'b10), .state({trees[1242], lumberyards[1242]}));
acre acre_24_43 (.clk(clk), .en(en), .top_left({trees[1192], lumberyards[1192]}), .top({trees[1193], lumberyards[1193]}), .top_right({trees[1194], lumberyards[1194]}), .left({trees[1242], lumberyards[1242]}), .right({trees[1244], lumberyards[1244]}), .bottom_left({trees[1292], lumberyards[1292]}), .bottom({trees[1293], lumberyards[1293]}), .bottom_right({trees[1294], lumberyards[1294]}), .init(2'b00), .state({trees[1243], lumberyards[1243]}));
acre acre_24_44 (.clk(clk), .en(en), .top_left({trees[1193], lumberyards[1193]}), .top({trees[1194], lumberyards[1194]}), .top_right({trees[1195], lumberyards[1195]}), .left({trees[1243], lumberyards[1243]}), .right({trees[1245], lumberyards[1245]}), .bottom_left({trees[1293], lumberyards[1293]}), .bottom({trees[1294], lumberyards[1294]}), .bottom_right({trees[1295], lumberyards[1295]}), .init(2'b00), .state({trees[1244], lumberyards[1244]}));
acre acre_24_45 (.clk(clk), .en(en), .top_left({trees[1194], lumberyards[1194]}), .top({trees[1195], lumberyards[1195]}), .top_right({trees[1196], lumberyards[1196]}), .left({trees[1244], lumberyards[1244]}), .right({trees[1246], lumberyards[1246]}), .bottom_left({trees[1294], lumberyards[1294]}), .bottom({trees[1295], lumberyards[1295]}), .bottom_right({trees[1296], lumberyards[1296]}), .init(2'b01), .state({trees[1245], lumberyards[1245]}));
acre acre_24_46 (.clk(clk), .en(en), .top_left({trees[1195], lumberyards[1195]}), .top({trees[1196], lumberyards[1196]}), .top_right({trees[1197], lumberyards[1197]}), .left({trees[1245], lumberyards[1245]}), .right({trees[1247], lumberyards[1247]}), .bottom_left({trees[1295], lumberyards[1295]}), .bottom({trees[1296], lumberyards[1296]}), .bottom_right({trees[1297], lumberyards[1297]}), .init(2'b00), .state({trees[1246], lumberyards[1246]}));
acre acre_24_47 (.clk(clk), .en(en), .top_left({trees[1196], lumberyards[1196]}), .top({trees[1197], lumberyards[1197]}), .top_right({trees[1198], lumberyards[1198]}), .left({trees[1246], lumberyards[1246]}), .right({trees[1248], lumberyards[1248]}), .bottom_left({trees[1296], lumberyards[1296]}), .bottom({trees[1297], lumberyards[1297]}), .bottom_right({trees[1298], lumberyards[1298]}), .init(2'b01), .state({trees[1247], lumberyards[1247]}));
acre acre_24_48 (.clk(clk), .en(en), .top_left({trees[1197], lumberyards[1197]}), .top({trees[1198], lumberyards[1198]}), .top_right({trees[1199], lumberyards[1199]}), .left({trees[1247], lumberyards[1247]}), .right({trees[1249], lumberyards[1249]}), .bottom_left({trees[1297], lumberyards[1297]}), .bottom({trees[1298], lumberyards[1298]}), .bottom_right({trees[1299], lumberyards[1299]}), .init(2'b10), .state({trees[1248], lumberyards[1248]}));
acre acre_24_49 (.clk(clk), .en(en), .top_left({trees[1198], lumberyards[1198]}), .top({trees[1199], lumberyards[1199]}), .top_right(2'b0), .left({trees[1248], lumberyards[1248]}), .right(2'b0), .bottom_left({trees[1298], lumberyards[1298]}), .bottom({trees[1299], lumberyards[1299]}), .bottom_right(2'b0), .init(2'b00), .state({trees[1249], lumberyards[1249]}));
acre acre_25_0 (.clk(clk), .en(en), .top_left(2'b0), .top({trees[1200], lumberyards[1200]}), .top_right({trees[1201], lumberyards[1201]}), .left(2'b0), .right({trees[1251], lumberyards[1251]}), .bottom_left(2'b0), .bottom({trees[1300], lumberyards[1300]}), .bottom_right({trees[1301], lumberyards[1301]}), .init(2'b10), .state({trees[1250], lumberyards[1250]}));
acre acre_25_1 (.clk(clk), .en(en), .top_left({trees[1200], lumberyards[1200]}), .top({trees[1201], lumberyards[1201]}), .top_right({trees[1202], lumberyards[1202]}), .left({trees[1250], lumberyards[1250]}), .right({trees[1252], lumberyards[1252]}), .bottom_left({trees[1300], lumberyards[1300]}), .bottom({trees[1301], lumberyards[1301]}), .bottom_right({trees[1302], lumberyards[1302]}), .init(2'b00), .state({trees[1251], lumberyards[1251]}));
acre acre_25_2 (.clk(clk), .en(en), .top_left({trees[1201], lumberyards[1201]}), .top({trees[1202], lumberyards[1202]}), .top_right({trees[1203], lumberyards[1203]}), .left({trees[1251], lumberyards[1251]}), .right({trees[1253], lumberyards[1253]}), .bottom_left({trees[1301], lumberyards[1301]}), .bottom({trees[1302], lumberyards[1302]}), .bottom_right({trees[1303], lumberyards[1303]}), .init(2'b00), .state({trees[1252], lumberyards[1252]}));
acre acre_25_3 (.clk(clk), .en(en), .top_left({trees[1202], lumberyards[1202]}), .top({trees[1203], lumberyards[1203]}), .top_right({trees[1204], lumberyards[1204]}), .left({trees[1252], lumberyards[1252]}), .right({trees[1254], lumberyards[1254]}), .bottom_left({trees[1302], lumberyards[1302]}), .bottom({trees[1303], lumberyards[1303]}), .bottom_right({trees[1304], lumberyards[1304]}), .init(2'b00), .state({trees[1253], lumberyards[1253]}));
acre acre_25_4 (.clk(clk), .en(en), .top_left({trees[1203], lumberyards[1203]}), .top({trees[1204], lumberyards[1204]}), .top_right({trees[1205], lumberyards[1205]}), .left({trees[1253], lumberyards[1253]}), .right({trees[1255], lumberyards[1255]}), .bottom_left({trees[1303], lumberyards[1303]}), .bottom({trees[1304], lumberyards[1304]}), .bottom_right({trees[1305], lumberyards[1305]}), .init(2'b00), .state({trees[1254], lumberyards[1254]}));
acre acre_25_5 (.clk(clk), .en(en), .top_left({trees[1204], lumberyards[1204]}), .top({trees[1205], lumberyards[1205]}), .top_right({trees[1206], lumberyards[1206]}), .left({trees[1254], lumberyards[1254]}), .right({trees[1256], lumberyards[1256]}), .bottom_left({trees[1304], lumberyards[1304]}), .bottom({trees[1305], lumberyards[1305]}), .bottom_right({trees[1306], lumberyards[1306]}), .init(2'b00), .state({trees[1255], lumberyards[1255]}));
acre acre_25_6 (.clk(clk), .en(en), .top_left({trees[1205], lumberyards[1205]}), .top({trees[1206], lumberyards[1206]}), .top_right({trees[1207], lumberyards[1207]}), .left({trees[1255], lumberyards[1255]}), .right({trees[1257], lumberyards[1257]}), .bottom_left({trees[1305], lumberyards[1305]}), .bottom({trees[1306], lumberyards[1306]}), .bottom_right({trees[1307], lumberyards[1307]}), .init(2'b01), .state({trees[1256], lumberyards[1256]}));
acre acre_25_7 (.clk(clk), .en(en), .top_left({trees[1206], lumberyards[1206]}), .top({trees[1207], lumberyards[1207]}), .top_right({trees[1208], lumberyards[1208]}), .left({trees[1256], lumberyards[1256]}), .right({trees[1258], lumberyards[1258]}), .bottom_left({trees[1306], lumberyards[1306]}), .bottom({trees[1307], lumberyards[1307]}), .bottom_right({trees[1308], lumberyards[1308]}), .init(2'b00), .state({trees[1257], lumberyards[1257]}));
acre acre_25_8 (.clk(clk), .en(en), .top_left({trees[1207], lumberyards[1207]}), .top({trees[1208], lumberyards[1208]}), .top_right({trees[1209], lumberyards[1209]}), .left({trees[1257], lumberyards[1257]}), .right({trees[1259], lumberyards[1259]}), .bottom_left({trees[1307], lumberyards[1307]}), .bottom({trees[1308], lumberyards[1308]}), .bottom_right({trees[1309], lumberyards[1309]}), .init(2'b00), .state({trees[1258], lumberyards[1258]}));
acre acre_25_9 (.clk(clk), .en(en), .top_left({trees[1208], lumberyards[1208]}), .top({trees[1209], lumberyards[1209]}), .top_right({trees[1210], lumberyards[1210]}), .left({trees[1258], lumberyards[1258]}), .right({trees[1260], lumberyards[1260]}), .bottom_left({trees[1308], lumberyards[1308]}), .bottom({trees[1309], lumberyards[1309]}), .bottom_right({trees[1310], lumberyards[1310]}), .init(2'b00), .state({trees[1259], lumberyards[1259]}));
acre acre_25_10 (.clk(clk), .en(en), .top_left({trees[1209], lumberyards[1209]}), .top({trees[1210], lumberyards[1210]}), .top_right({trees[1211], lumberyards[1211]}), .left({trees[1259], lumberyards[1259]}), .right({trees[1261], lumberyards[1261]}), .bottom_left({trees[1309], lumberyards[1309]}), .bottom({trees[1310], lumberyards[1310]}), .bottom_right({trees[1311], lumberyards[1311]}), .init(2'b01), .state({trees[1260], lumberyards[1260]}));
acre acre_25_11 (.clk(clk), .en(en), .top_left({trees[1210], lumberyards[1210]}), .top({trees[1211], lumberyards[1211]}), .top_right({trees[1212], lumberyards[1212]}), .left({trees[1260], lumberyards[1260]}), .right({trees[1262], lumberyards[1262]}), .bottom_left({trees[1310], lumberyards[1310]}), .bottom({trees[1311], lumberyards[1311]}), .bottom_right({trees[1312], lumberyards[1312]}), .init(2'b01), .state({trees[1261], lumberyards[1261]}));
acre acre_25_12 (.clk(clk), .en(en), .top_left({trees[1211], lumberyards[1211]}), .top({trees[1212], lumberyards[1212]}), .top_right({trees[1213], lumberyards[1213]}), .left({trees[1261], lumberyards[1261]}), .right({trees[1263], lumberyards[1263]}), .bottom_left({trees[1311], lumberyards[1311]}), .bottom({trees[1312], lumberyards[1312]}), .bottom_right({trees[1313], lumberyards[1313]}), .init(2'b00), .state({trees[1262], lumberyards[1262]}));
acre acre_25_13 (.clk(clk), .en(en), .top_left({trees[1212], lumberyards[1212]}), .top({trees[1213], lumberyards[1213]}), .top_right({trees[1214], lumberyards[1214]}), .left({trees[1262], lumberyards[1262]}), .right({trees[1264], lumberyards[1264]}), .bottom_left({trees[1312], lumberyards[1312]}), .bottom({trees[1313], lumberyards[1313]}), .bottom_right({trees[1314], lumberyards[1314]}), .init(2'b00), .state({trees[1263], lumberyards[1263]}));
acre acre_25_14 (.clk(clk), .en(en), .top_left({trees[1213], lumberyards[1213]}), .top({trees[1214], lumberyards[1214]}), .top_right({trees[1215], lumberyards[1215]}), .left({trees[1263], lumberyards[1263]}), .right({trees[1265], lumberyards[1265]}), .bottom_left({trees[1313], lumberyards[1313]}), .bottom({trees[1314], lumberyards[1314]}), .bottom_right({trees[1315], lumberyards[1315]}), .init(2'b00), .state({trees[1264], lumberyards[1264]}));
acre acre_25_15 (.clk(clk), .en(en), .top_left({trees[1214], lumberyards[1214]}), .top({trees[1215], lumberyards[1215]}), .top_right({trees[1216], lumberyards[1216]}), .left({trees[1264], lumberyards[1264]}), .right({trees[1266], lumberyards[1266]}), .bottom_left({trees[1314], lumberyards[1314]}), .bottom({trees[1315], lumberyards[1315]}), .bottom_right({trees[1316], lumberyards[1316]}), .init(2'b00), .state({trees[1265], lumberyards[1265]}));
acre acre_25_16 (.clk(clk), .en(en), .top_left({trees[1215], lumberyards[1215]}), .top({trees[1216], lumberyards[1216]}), .top_right({trees[1217], lumberyards[1217]}), .left({trees[1265], lumberyards[1265]}), .right({trees[1267], lumberyards[1267]}), .bottom_left({trees[1315], lumberyards[1315]}), .bottom({trees[1316], lumberyards[1316]}), .bottom_right({trees[1317], lumberyards[1317]}), .init(2'b00), .state({trees[1266], lumberyards[1266]}));
acre acre_25_17 (.clk(clk), .en(en), .top_left({trees[1216], lumberyards[1216]}), .top({trees[1217], lumberyards[1217]}), .top_right({trees[1218], lumberyards[1218]}), .left({trees[1266], lumberyards[1266]}), .right({trees[1268], lumberyards[1268]}), .bottom_left({trees[1316], lumberyards[1316]}), .bottom({trees[1317], lumberyards[1317]}), .bottom_right({trees[1318], lumberyards[1318]}), .init(2'b10), .state({trees[1267], lumberyards[1267]}));
acre acre_25_18 (.clk(clk), .en(en), .top_left({trees[1217], lumberyards[1217]}), .top({trees[1218], lumberyards[1218]}), .top_right({trees[1219], lumberyards[1219]}), .left({trees[1267], lumberyards[1267]}), .right({trees[1269], lumberyards[1269]}), .bottom_left({trees[1317], lumberyards[1317]}), .bottom({trees[1318], lumberyards[1318]}), .bottom_right({trees[1319], lumberyards[1319]}), .init(2'b00), .state({trees[1268], lumberyards[1268]}));
acre acre_25_19 (.clk(clk), .en(en), .top_left({trees[1218], lumberyards[1218]}), .top({trees[1219], lumberyards[1219]}), .top_right({trees[1220], lumberyards[1220]}), .left({trees[1268], lumberyards[1268]}), .right({trees[1270], lumberyards[1270]}), .bottom_left({trees[1318], lumberyards[1318]}), .bottom({trees[1319], lumberyards[1319]}), .bottom_right({trees[1320], lumberyards[1320]}), .init(2'b00), .state({trees[1269], lumberyards[1269]}));
acre acre_25_20 (.clk(clk), .en(en), .top_left({trees[1219], lumberyards[1219]}), .top({trees[1220], lumberyards[1220]}), .top_right({trees[1221], lumberyards[1221]}), .left({trees[1269], lumberyards[1269]}), .right({trees[1271], lumberyards[1271]}), .bottom_left({trees[1319], lumberyards[1319]}), .bottom({trees[1320], lumberyards[1320]}), .bottom_right({trees[1321], lumberyards[1321]}), .init(2'b10), .state({trees[1270], lumberyards[1270]}));
acre acre_25_21 (.clk(clk), .en(en), .top_left({trees[1220], lumberyards[1220]}), .top({trees[1221], lumberyards[1221]}), .top_right({trees[1222], lumberyards[1222]}), .left({trees[1270], lumberyards[1270]}), .right({trees[1272], lumberyards[1272]}), .bottom_left({trees[1320], lumberyards[1320]}), .bottom({trees[1321], lumberyards[1321]}), .bottom_right({trees[1322], lumberyards[1322]}), .init(2'b00), .state({trees[1271], lumberyards[1271]}));
acre acre_25_22 (.clk(clk), .en(en), .top_left({trees[1221], lumberyards[1221]}), .top({trees[1222], lumberyards[1222]}), .top_right({trees[1223], lumberyards[1223]}), .left({trees[1271], lumberyards[1271]}), .right({trees[1273], lumberyards[1273]}), .bottom_left({trees[1321], lumberyards[1321]}), .bottom({trees[1322], lumberyards[1322]}), .bottom_right({trees[1323], lumberyards[1323]}), .init(2'b00), .state({trees[1272], lumberyards[1272]}));
acre acre_25_23 (.clk(clk), .en(en), .top_left({trees[1222], lumberyards[1222]}), .top({trees[1223], lumberyards[1223]}), .top_right({trees[1224], lumberyards[1224]}), .left({trees[1272], lumberyards[1272]}), .right({trees[1274], lumberyards[1274]}), .bottom_left({trees[1322], lumberyards[1322]}), .bottom({trees[1323], lumberyards[1323]}), .bottom_right({trees[1324], lumberyards[1324]}), .init(2'b00), .state({trees[1273], lumberyards[1273]}));
acre acre_25_24 (.clk(clk), .en(en), .top_left({trees[1223], lumberyards[1223]}), .top({trees[1224], lumberyards[1224]}), .top_right({trees[1225], lumberyards[1225]}), .left({trees[1273], lumberyards[1273]}), .right({trees[1275], lumberyards[1275]}), .bottom_left({trees[1323], lumberyards[1323]}), .bottom({trees[1324], lumberyards[1324]}), .bottom_right({trees[1325], lumberyards[1325]}), .init(2'b01), .state({trees[1274], lumberyards[1274]}));
acre acre_25_25 (.clk(clk), .en(en), .top_left({trees[1224], lumberyards[1224]}), .top({trees[1225], lumberyards[1225]}), .top_right({trees[1226], lumberyards[1226]}), .left({trees[1274], lumberyards[1274]}), .right({trees[1276], lumberyards[1276]}), .bottom_left({trees[1324], lumberyards[1324]}), .bottom({trees[1325], lumberyards[1325]}), .bottom_right({trees[1326], lumberyards[1326]}), .init(2'b10), .state({trees[1275], lumberyards[1275]}));
acre acre_25_26 (.clk(clk), .en(en), .top_left({trees[1225], lumberyards[1225]}), .top({trees[1226], lumberyards[1226]}), .top_right({trees[1227], lumberyards[1227]}), .left({trees[1275], lumberyards[1275]}), .right({trees[1277], lumberyards[1277]}), .bottom_left({trees[1325], lumberyards[1325]}), .bottom({trees[1326], lumberyards[1326]}), .bottom_right({trees[1327], lumberyards[1327]}), .init(2'b01), .state({trees[1276], lumberyards[1276]}));
acre acre_25_27 (.clk(clk), .en(en), .top_left({trees[1226], lumberyards[1226]}), .top({trees[1227], lumberyards[1227]}), .top_right({trees[1228], lumberyards[1228]}), .left({trees[1276], lumberyards[1276]}), .right({trees[1278], lumberyards[1278]}), .bottom_left({trees[1326], lumberyards[1326]}), .bottom({trees[1327], lumberyards[1327]}), .bottom_right({trees[1328], lumberyards[1328]}), .init(2'b00), .state({trees[1277], lumberyards[1277]}));
acre acre_25_28 (.clk(clk), .en(en), .top_left({trees[1227], lumberyards[1227]}), .top({trees[1228], lumberyards[1228]}), .top_right({trees[1229], lumberyards[1229]}), .left({trees[1277], lumberyards[1277]}), .right({trees[1279], lumberyards[1279]}), .bottom_left({trees[1327], lumberyards[1327]}), .bottom({trees[1328], lumberyards[1328]}), .bottom_right({trees[1329], lumberyards[1329]}), .init(2'b01), .state({trees[1278], lumberyards[1278]}));
acre acre_25_29 (.clk(clk), .en(en), .top_left({trees[1228], lumberyards[1228]}), .top({trees[1229], lumberyards[1229]}), .top_right({trees[1230], lumberyards[1230]}), .left({trees[1278], lumberyards[1278]}), .right({trees[1280], lumberyards[1280]}), .bottom_left({trees[1328], lumberyards[1328]}), .bottom({trees[1329], lumberyards[1329]}), .bottom_right({trees[1330], lumberyards[1330]}), .init(2'b00), .state({trees[1279], lumberyards[1279]}));
acre acre_25_30 (.clk(clk), .en(en), .top_left({trees[1229], lumberyards[1229]}), .top({trees[1230], lumberyards[1230]}), .top_right({trees[1231], lumberyards[1231]}), .left({trees[1279], lumberyards[1279]}), .right({trees[1281], lumberyards[1281]}), .bottom_left({trees[1329], lumberyards[1329]}), .bottom({trees[1330], lumberyards[1330]}), .bottom_right({trees[1331], lumberyards[1331]}), .init(2'b00), .state({trees[1280], lumberyards[1280]}));
acre acre_25_31 (.clk(clk), .en(en), .top_left({trees[1230], lumberyards[1230]}), .top({trees[1231], lumberyards[1231]}), .top_right({trees[1232], lumberyards[1232]}), .left({trees[1280], lumberyards[1280]}), .right({trees[1282], lumberyards[1282]}), .bottom_left({trees[1330], lumberyards[1330]}), .bottom({trees[1331], lumberyards[1331]}), .bottom_right({trees[1332], lumberyards[1332]}), .init(2'b00), .state({trees[1281], lumberyards[1281]}));
acre acre_25_32 (.clk(clk), .en(en), .top_left({trees[1231], lumberyards[1231]}), .top({trees[1232], lumberyards[1232]}), .top_right({trees[1233], lumberyards[1233]}), .left({trees[1281], lumberyards[1281]}), .right({trees[1283], lumberyards[1283]}), .bottom_left({trees[1331], lumberyards[1331]}), .bottom({trees[1332], lumberyards[1332]}), .bottom_right({trees[1333], lumberyards[1333]}), .init(2'b00), .state({trees[1282], lumberyards[1282]}));
acre acre_25_33 (.clk(clk), .en(en), .top_left({trees[1232], lumberyards[1232]}), .top({trees[1233], lumberyards[1233]}), .top_right({trees[1234], lumberyards[1234]}), .left({trees[1282], lumberyards[1282]}), .right({trees[1284], lumberyards[1284]}), .bottom_left({trees[1332], lumberyards[1332]}), .bottom({trees[1333], lumberyards[1333]}), .bottom_right({trees[1334], lumberyards[1334]}), .init(2'b10), .state({trees[1283], lumberyards[1283]}));
acre acre_25_34 (.clk(clk), .en(en), .top_left({trees[1233], lumberyards[1233]}), .top({trees[1234], lumberyards[1234]}), .top_right({trees[1235], lumberyards[1235]}), .left({trees[1283], lumberyards[1283]}), .right({trees[1285], lumberyards[1285]}), .bottom_left({trees[1333], lumberyards[1333]}), .bottom({trees[1334], lumberyards[1334]}), .bottom_right({trees[1335], lumberyards[1335]}), .init(2'b01), .state({trees[1284], lumberyards[1284]}));
acre acre_25_35 (.clk(clk), .en(en), .top_left({trees[1234], lumberyards[1234]}), .top({trees[1235], lumberyards[1235]}), .top_right({trees[1236], lumberyards[1236]}), .left({trees[1284], lumberyards[1284]}), .right({trees[1286], lumberyards[1286]}), .bottom_left({trees[1334], lumberyards[1334]}), .bottom({trees[1335], lumberyards[1335]}), .bottom_right({trees[1336], lumberyards[1336]}), .init(2'b00), .state({trees[1285], lumberyards[1285]}));
acre acre_25_36 (.clk(clk), .en(en), .top_left({trees[1235], lumberyards[1235]}), .top({trees[1236], lumberyards[1236]}), .top_right({trees[1237], lumberyards[1237]}), .left({trees[1285], lumberyards[1285]}), .right({trees[1287], lumberyards[1287]}), .bottom_left({trees[1335], lumberyards[1335]}), .bottom({trees[1336], lumberyards[1336]}), .bottom_right({trees[1337], lumberyards[1337]}), .init(2'b00), .state({trees[1286], lumberyards[1286]}));
acre acre_25_37 (.clk(clk), .en(en), .top_left({trees[1236], lumberyards[1236]}), .top({trees[1237], lumberyards[1237]}), .top_right({trees[1238], lumberyards[1238]}), .left({trees[1286], lumberyards[1286]}), .right({trees[1288], lumberyards[1288]}), .bottom_left({trees[1336], lumberyards[1336]}), .bottom({trees[1337], lumberyards[1337]}), .bottom_right({trees[1338], lumberyards[1338]}), .init(2'b10), .state({trees[1287], lumberyards[1287]}));
acre acre_25_38 (.clk(clk), .en(en), .top_left({trees[1237], lumberyards[1237]}), .top({trees[1238], lumberyards[1238]}), .top_right({trees[1239], lumberyards[1239]}), .left({trees[1287], lumberyards[1287]}), .right({trees[1289], lumberyards[1289]}), .bottom_left({trees[1337], lumberyards[1337]}), .bottom({trees[1338], lumberyards[1338]}), .bottom_right({trees[1339], lumberyards[1339]}), .init(2'b01), .state({trees[1288], lumberyards[1288]}));
acre acre_25_39 (.clk(clk), .en(en), .top_left({trees[1238], lumberyards[1238]}), .top({trees[1239], lumberyards[1239]}), .top_right({trees[1240], lumberyards[1240]}), .left({trees[1288], lumberyards[1288]}), .right({trees[1290], lumberyards[1290]}), .bottom_left({trees[1338], lumberyards[1338]}), .bottom({trees[1339], lumberyards[1339]}), .bottom_right({trees[1340], lumberyards[1340]}), .init(2'b00), .state({trees[1289], lumberyards[1289]}));
acre acre_25_40 (.clk(clk), .en(en), .top_left({trees[1239], lumberyards[1239]}), .top({trees[1240], lumberyards[1240]}), .top_right({trees[1241], lumberyards[1241]}), .left({trees[1289], lumberyards[1289]}), .right({trees[1291], lumberyards[1291]}), .bottom_left({trees[1339], lumberyards[1339]}), .bottom({trees[1340], lumberyards[1340]}), .bottom_right({trees[1341], lumberyards[1341]}), .init(2'b00), .state({trees[1290], lumberyards[1290]}));
acre acre_25_41 (.clk(clk), .en(en), .top_left({trees[1240], lumberyards[1240]}), .top({trees[1241], lumberyards[1241]}), .top_right({trees[1242], lumberyards[1242]}), .left({trees[1290], lumberyards[1290]}), .right({trees[1292], lumberyards[1292]}), .bottom_left({trees[1340], lumberyards[1340]}), .bottom({trees[1341], lumberyards[1341]}), .bottom_right({trees[1342], lumberyards[1342]}), .init(2'b00), .state({trees[1291], lumberyards[1291]}));
acre acre_25_42 (.clk(clk), .en(en), .top_left({trees[1241], lumberyards[1241]}), .top({trees[1242], lumberyards[1242]}), .top_right({trees[1243], lumberyards[1243]}), .left({trees[1291], lumberyards[1291]}), .right({trees[1293], lumberyards[1293]}), .bottom_left({trees[1341], lumberyards[1341]}), .bottom({trees[1342], lumberyards[1342]}), .bottom_right({trees[1343], lumberyards[1343]}), .init(2'b10), .state({trees[1292], lumberyards[1292]}));
acre acre_25_43 (.clk(clk), .en(en), .top_left({trees[1242], lumberyards[1242]}), .top({trees[1243], lumberyards[1243]}), .top_right({trees[1244], lumberyards[1244]}), .left({trees[1292], lumberyards[1292]}), .right({trees[1294], lumberyards[1294]}), .bottom_left({trees[1342], lumberyards[1342]}), .bottom({trees[1343], lumberyards[1343]}), .bottom_right({trees[1344], lumberyards[1344]}), .init(2'b00), .state({trees[1293], lumberyards[1293]}));
acre acre_25_44 (.clk(clk), .en(en), .top_left({trees[1243], lumberyards[1243]}), .top({trees[1244], lumberyards[1244]}), .top_right({trees[1245], lumberyards[1245]}), .left({trees[1293], lumberyards[1293]}), .right({trees[1295], lumberyards[1295]}), .bottom_left({trees[1343], lumberyards[1343]}), .bottom({trees[1344], lumberyards[1344]}), .bottom_right({trees[1345], lumberyards[1345]}), .init(2'b00), .state({trees[1294], lumberyards[1294]}));
acre acre_25_45 (.clk(clk), .en(en), .top_left({trees[1244], lumberyards[1244]}), .top({trees[1245], lumberyards[1245]}), .top_right({trees[1246], lumberyards[1246]}), .left({trees[1294], lumberyards[1294]}), .right({trees[1296], lumberyards[1296]}), .bottom_left({trees[1344], lumberyards[1344]}), .bottom({trees[1345], lumberyards[1345]}), .bottom_right({trees[1346], lumberyards[1346]}), .init(2'b00), .state({trees[1295], lumberyards[1295]}));
acre acre_25_46 (.clk(clk), .en(en), .top_left({trees[1245], lumberyards[1245]}), .top({trees[1246], lumberyards[1246]}), .top_right({trees[1247], lumberyards[1247]}), .left({trees[1295], lumberyards[1295]}), .right({trees[1297], lumberyards[1297]}), .bottom_left({trees[1345], lumberyards[1345]}), .bottom({trees[1346], lumberyards[1346]}), .bottom_right({trees[1347], lumberyards[1347]}), .init(2'b00), .state({trees[1296], lumberyards[1296]}));
acre acre_25_47 (.clk(clk), .en(en), .top_left({trees[1246], lumberyards[1246]}), .top({trees[1247], lumberyards[1247]}), .top_right({trees[1248], lumberyards[1248]}), .left({trees[1296], lumberyards[1296]}), .right({trees[1298], lumberyards[1298]}), .bottom_left({trees[1346], lumberyards[1346]}), .bottom({trees[1347], lumberyards[1347]}), .bottom_right({trees[1348], lumberyards[1348]}), .init(2'b10), .state({trees[1297], lumberyards[1297]}));
acre acre_25_48 (.clk(clk), .en(en), .top_left({trees[1247], lumberyards[1247]}), .top({trees[1248], lumberyards[1248]}), .top_right({trees[1249], lumberyards[1249]}), .left({trees[1297], lumberyards[1297]}), .right({trees[1299], lumberyards[1299]}), .bottom_left({trees[1347], lumberyards[1347]}), .bottom({trees[1348], lumberyards[1348]}), .bottom_right({trees[1349], lumberyards[1349]}), .init(2'b00), .state({trees[1298], lumberyards[1298]}));
acre acre_25_49 (.clk(clk), .en(en), .top_left({trees[1248], lumberyards[1248]}), .top({trees[1249], lumberyards[1249]}), .top_right(2'b0), .left({trees[1298], lumberyards[1298]}), .right(2'b0), .bottom_left({trees[1348], lumberyards[1348]}), .bottom({trees[1349], lumberyards[1349]}), .bottom_right(2'b0), .init(2'b00), .state({trees[1299], lumberyards[1299]}));
acre acre_26_0 (.clk(clk), .en(en), .top_left(2'b0), .top({trees[1250], lumberyards[1250]}), .top_right({trees[1251], lumberyards[1251]}), .left(2'b0), .right({trees[1301], lumberyards[1301]}), .bottom_left(2'b0), .bottom({trees[1350], lumberyards[1350]}), .bottom_right({trees[1351], lumberyards[1351]}), .init(2'b10), .state({trees[1300], lumberyards[1300]}));
acre acre_26_1 (.clk(clk), .en(en), .top_left({trees[1250], lumberyards[1250]}), .top({trees[1251], lumberyards[1251]}), .top_right({trees[1252], lumberyards[1252]}), .left({trees[1300], lumberyards[1300]}), .right({trees[1302], lumberyards[1302]}), .bottom_left({trees[1350], lumberyards[1350]}), .bottom({trees[1351], lumberyards[1351]}), .bottom_right({trees[1352], lumberyards[1352]}), .init(2'b00), .state({trees[1301], lumberyards[1301]}));
acre acre_26_2 (.clk(clk), .en(en), .top_left({trees[1251], lumberyards[1251]}), .top({trees[1252], lumberyards[1252]}), .top_right({trees[1253], lumberyards[1253]}), .left({trees[1301], lumberyards[1301]}), .right({trees[1303], lumberyards[1303]}), .bottom_left({trees[1351], lumberyards[1351]}), .bottom({trees[1352], lumberyards[1352]}), .bottom_right({trees[1353], lumberyards[1353]}), .init(2'b00), .state({trees[1302], lumberyards[1302]}));
acre acre_26_3 (.clk(clk), .en(en), .top_left({trees[1252], lumberyards[1252]}), .top({trees[1253], lumberyards[1253]}), .top_right({trees[1254], lumberyards[1254]}), .left({trees[1302], lumberyards[1302]}), .right({trees[1304], lumberyards[1304]}), .bottom_left({trees[1352], lumberyards[1352]}), .bottom({trees[1353], lumberyards[1353]}), .bottom_right({trees[1354], lumberyards[1354]}), .init(2'b10), .state({trees[1303], lumberyards[1303]}));
acre acre_26_4 (.clk(clk), .en(en), .top_left({trees[1253], lumberyards[1253]}), .top({trees[1254], lumberyards[1254]}), .top_right({trees[1255], lumberyards[1255]}), .left({trees[1303], lumberyards[1303]}), .right({trees[1305], lumberyards[1305]}), .bottom_left({trees[1353], lumberyards[1353]}), .bottom({trees[1354], lumberyards[1354]}), .bottom_right({trees[1355], lumberyards[1355]}), .init(2'b00), .state({trees[1304], lumberyards[1304]}));
acre acre_26_5 (.clk(clk), .en(en), .top_left({trees[1254], lumberyards[1254]}), .top({trees[1255], lumberyards[1255]}), .top_right({trees[1256], lumberyards[1256]}), .left({trees[1304], lumberyards[1304]}), .right({trees[1306], lumberyards[1306]}), .bottom_left({trees[1354], lumberyards[1354]}), .bottom({trees[1355], lumberyards[1355]}), .bottom_right({trees[1356], lumberyards[1356]}), .init(2'b00), .state({trees[1305], lumberyards[1305]}));
acre acre_26_6 (.clk(clk), .en(en), .top_left({trees[1255], lumberyards[1255]}), .top({trees[1256], lumberyards[1256]}), .top_right({trees[1257], lumberyards[1257]}), .left({trees[1305], lumberyards[1305]}), .right({trees[1307], lumberyards[1307]}), .bottom_left({trees[1355], lumberyards[1355]}), .bottom({trees[1356], lumberyards[1356]}), .bottom_right({trees[1357], lumberyards[1357]}), .init(2'b00), .state({trees[1306], lumberyards[1306]}));
acre acre_26_7 (.clk(clk), .en(en), .top_left({trees[1256], lumberyards[1256]}), .top({trees[1257], lumberyards[1257]}), .top_right({trees[1258], lumberyards[1258]}), .left({trees[1306], lumberyards[1306]}), .right({trees[1308], lumberyards[1308]}), .bottom_left({trees[1356], lumberyards[1356]}), .bottom({trees[1357], lumberyards[1357]}), .bottom_right({trees[1358], lumberyards[1358]}), .init(2'b00), .state({trees[1307], lumberyards[1307]}));
acre acre_26_8 (.clk(clk), .en(en), .top_left({trees[1257], lumberyards[1257]}), .top({trees[1258], lumberyards[1258]}), .top_right({trees[1259], lumberyards[1259]}), .left({trees[1307], lumberyards[1307]}), .right({trees[1309], lumberyards[1309]}), .bottom_left({trees[1357], lumberyards[1357]}), .bottom({trees[1358], lumberyards[1358]}), .bottom_right({trees[1359], lumberyards[1359]}), .init(2'b10), .state({trees[1308], lumberyards[1308]}));
acre acre_26_9 (.clk(clk), .en(en), .top_left({trees[1258], lumberyards[1258]}), .top({trees[1259], lumberyards[1259]}), .top_right({trees[1260], lumberyards[1260]}), .left({trees[1308], lumberyards[1308]}), .right({trees[1310], lumberyards[1310]}), .bottom_left({trees[1358], lumberyards[1358]}), .bottom({trees[1359], lumberyards[1359]}), .bottom_right({trees[1360], lumberyards[1360]}), .init(2'b00), .state({trees[1309], lumberyards[1309]}));
acre acre_26_10 (.clk(clk), .en(en), .top_left({trees[1259], lumberyards[1259]}), .top({trees[1260], lumberyards[1260]}), .top_right({trees[1261], lumberyards[1261]}), .left({trees[1309], lumberyards[1309]}), .right({trees[1311], lumberyards[1311]}), .bottom_left({trees[1359], lumberyards[1359]}), .bottom({trees[1360], lumberyards[1360]}), .bottom_right({trees[1361], lumberyards[1361]}), .init(2'b00), .state({trees[1310], lumberyards[1310]}));
acre acre_26_11 (.clk(clk), .en(en), .top_left({trees[1260], lumberyards[1260]}), .top({trees[1261], lumberyards[1261]}), .top_right({trees[1262], lumberyards[1262]}), .left({trees[1310], lumberyards[1310]}), .right({trees[1312], lumberyards[1312]}), .bottom_left({trees[1360], lumberyards[1360]}), .bottom({trees[1361], lumberyards[1361]}), .bottom_right({trees[1362], lumberyards[1362]}), .init(2'b00), .state({trees[1311], lumberyards[1311]}));
acre acre_26_12 (.clk(clk), .en(en), .top_left({trees[1261], lumberyards[1261]}), .top({trees[1262], lumberyards[1262]}), .top_right({trees[1263], lumberyards[1263]}), .left({trees[1311], lumberyards[1311]}), .right({trees[1313], lumberyards[1313]}), .bottom_left({trees[1361], lumberyards[1361]}), .bottom({trees[1362], lumberyards[1362]}), .bottom_right({trees[1363], lumberyards[1363]}), .init(2'b01), .state({trees[1312], lumberyards[1312]}));
acre acre_26_13 (.clk(clk), .en(en), .top_left({trees[1262], lumberyards[1262]}), .top({trees[1263], lumberyards[1263]}), .top_right({trees[1264], lumberyards[1264]}), .left({trees[1312], lumberyards[1312]}), .right({trees[1314], lumberyards[1314]}), .bottom_left({trees[1362], lumberyards[1362]}), .bottom({trees[1363], lumberyards[1363]}), .bottom_right({trees[1364], lumberyards[1364]}), .init(2'b01), .state({trees[1313], lumberyards[1313]}));
acre acre_26_14 (.clk(clk), .en(en), .top_left({trees[1263], lumberyards[1263]}), .top({trees[1264], lumberyards[1264]}), .top_right({trees[1265], lumberyards[1265]}), .left({trees[1313], lumberyards[1313]}), .right({trees[1315], lumberyards[1315]}), .bottom_left({trees[1363], lumberyards[1363]}), .bottom({trees[1364], lumberyards[1364]}), .bottom_right({trees[1365], lumberyards[1365]}), .init(2'b00), .state({trees[1314], lumberyards[1314]}));
acre acre_26_15 (.clk(clk), .en(en), .top_left({trees[1264], lumberyards[1264]}), .top({trees[1265], lumberyards[1265]}), .top_right({trees[1266], lumberyards[1266]}), .left({trees[1314], lumberyards[1314]}), .right({trees[1316], lumberyards[1316]}), .bottom_left({trees[1364], lumberyards[1364]}), .bottom({trees[1365], lumberyards[1365]}), .bottom_right({trees[1366], lumberyards[1366]}), .init(2'b10), .state({trees[1315], lumberyards[1315]}));
acre acre_26_16 (.clk(clk), .en(en), .top_left({trees[1265], lumberyards[1265]}), .top({trees[1266], lumberyards[1266]}), .top_right({trees[1267], lumberyards[1267]}), .left({trees[1315], lumberyards[1315]}), .right({trees[1317], lumberyards[1317]}), .bottom_left({trees[1365], lumberyards[1365]}), .bottom({trees[1366], lumberyards[1366]}), .bottom_right({trees[1367], lumberyards[1367]}), .init(2'b00), .state({trees[1316], lumberyards[1316]}));
acre acre_26_17 (.clk(clk), .en(en), .top_left({trees[1266], lumberyards[1266]}), .top({trees[1267], lumberyards[1267]}), .top_right({trees[1268], lumberyards[1268]}), .left({trees[1316], lumberyards[1316]}), .right({trees[1318], lumberyards[1318]}), .bottom_left({trees[1366], lumberyards[1366]}), .bottom({trees[1367], lumberyards[1367]}), .bottom_right({trees[1368], lumberyards[1368]}), .init(2'b00), .state({trees[1317], lumberyards[1317]}));
acre acre_26_18 (.clk(clk), .en(en), .top_left({trees[1267], lumberyards[1267]}), .top({trees[1268], lumberyards[1268]}), .top_right({trees[1269], lumberyards[1269]}), .left({trees[1317], lumberyards[1317]}), .right({trees[1319], lumberyards[1319]}), .bottom_left({trees[1367], lumberyards[1367]}), .bottom({trees[1368], lumberyards[1368]}), .bottom_right({trees[1369], lumberyards[1369]}), .init(2'b00), .state({trees[1318], lumberyards[1318]}));
acre acre_26_19 (.clk(clk), .en(en), .top_left({trees[1268], lumberyards[1268]}), .top({trees[1269], lumberyards[1269]}), .top_right({trees[1270], lumberyards[1270]}), .left({trees[1318], lumberyards[1318]}), .right({trees[1320], lumberyards[1320]}), .bottom_left({trees[1368], lumberyards[1368]}), .bottom({trees[1369], lumberyards[1369]}), .bottom_right({trees[1370], lumberyards[1370]}), .init(2'b00), .state({trees[1319], lumberyards[1319]}));
acre acre_26_20 (.clk(clk), .en(en), .top_left({trees[1269], lumberyards[1269]}), .top({trees[1270], lumberyards[1270]}), .top_right({trees[1271], lumberyards[1271]}), .left({trees[1319], lumberyards[1319]}), .right({trees[1321], lumberyards[1321]}), .bottom_left({trees[1369], lumberyards[1369]}), .bottom({trees[1370], lumberyards[1370]}), .bottom_right({trees[1371], lumberyards[1371]}), .init(2'b00), .state({trees[1320], lumberyards[1320]}));
acre acre_26_21 (.clk(clk), .en(en), .top_left({trees[1270], lumberyards[1270]}), .top({trees[1271], lumberyards[1271]}), .top_right({trees[1272], lumberyards[1272]}), .left({trees[1320], lumberyards[1320]}), .right({trees[1322], lumberyards[1322]}), .bottom_left({trees[1370], lumberyards[1370]}), .bottom({trees[1371], lumberyards[1371]}), .bottom_right({trees[1372], lumberyards[1372]}), .init(2'b01), .state({trees[1321], lumberyards[1321]}));
acre acre_26_22 (.clk(clk), .en(en), .top_left({trees[1271], lumberyards[1271]}), .top({trees[1272], lumberyards[1272]}), .top_right({trees[1273], lumberyards[1273]}), .left({trees[1321], lumberyards[1321]}), .right({trees[1323], lumberyards[1323]}), .bottom_left({trees[1371], lumberyards[1371]}), .bottom({trees[1372], lumberyards[1372]}), .bottom_right({trees[1373], lumberyards[1373]}), .init(2'b10), .state({trees[1322], lumberyards[1322]}));
acre acre_26_23 (.clk(clk), .en(en), .top_left({trees[1272], lumberyards[1272]}), .top({trees[1273], lumberyards[1273]}), .top_right({trees[1274], lumberyards[1274]}), .left({trees[1322], lumberyards[1322]}), .right({trees[1324], lumberyards[1324]}), .bottom_left({trees[1372], lumberyards[1372]}), .bottom({trees[1373], lumberyards[1373]}), .bottom_right({trees[1374], lumberyards[1374]}), .init(2'b00), .state({trees[1323], lumberyards[1323]}));
acre acre_26_24 (.clk(clk), .en(en), .top_left({trees[1273], lumberyards[1273]}), .top({trees[1274], lumberyards[1274]}), .top_right({trees[1275], lumberyards[1275]}), .left({trees[1323], lumberyards[1323]}), .right({trees[1325], lumberyards[1325]}), .bottom_left({trees[1373], lumberyards[1373]}), .bottom({trees[1374], lumberyards[1374]}), .bottom_right({trees[1375], lumberyards[1375]}), .init(2'b01), .state({trees[1324], lumberyards[1324]}));
acre acre_26_25 (.clk(clk), .en(en), .top_left({trees[1274], lumberyards[1274]}), .top({trees[1275], lumberyards[1275]}), .top_right({trees[1276], lumberyards[1276]}), .left({trees[1324], lumberyards[1324]}), .right({trees[1326], lumberyards[1326]}), .bottom_left({trees[1374], lumberyards[1374]}), .bottom({trees[1375], lumberyards[1375]}), .bottom_right({trees[1376], lumberyards[1376]}), .init(2'b10), .state({trees[1325], lumberyards[1325]}));
acre acre_26_26 (.clk(clk), .en(en), .top_left({trees[1275], lumberyards[1275]}), .top({trees[1276], lumberyards[1276]}), .top_right({trees[1277], lumberyards[1277]}), .left({trees[1325], lumberyards[1325]}), .right({trees[1327], lumberyards[1327]}), .bottom_left({trees[1375], lumberyards[1375]}), .bottom({trees[1376], lumberyards[1376]}), .bottom_right({trees[1377], lumberyards[1377]}), .init(2'b00), .state({trees[1326], lumberyards[1326]}));
acre acre_26_27 (.clk(clk), .en(en), .top_left({trees[1276], lumberyards[1276]}), .top({trees[1277], lumberyards[1277]}), .top_right({trees[1278], lumberyards[1278]}), .left({trees[1326], lumberyards[1326]}), .right({trees[1328], lumberyards[1328]}), .bottom_left({trees[1376], lumberyards[1376]}), .bottom({trees[1377], lumberyards[1377]}), .bottom_right({trees[1378], lumberyards[1378]}), .init(2'b10), .state({trees[1327], lumberyards[1327]}));
acre acre_26_28 (.clk(clk), .en(en), .top_left({trees[1277], lumberyards[1277]}), .top({trees[1278], lumberyards[1278]}), .top_right({trees[1279], lumberyards[1279]}), .left({trees[1327], lumberyards[1327]}), .right({trees[1329], lumberyards[1329]}), .bottom_left({trees[1377], lumberyards[1377]}), .bottom({trees[1378], lumberyards[1378]}), .bottom_right({trees[1379], lumberyards[1379]}), .init(2'b10), .state({trees[1328], lumberyards[1328]}));
acre acre_26_29 (.clk(clk), .en(en), .top_left({trees[1278], lumberyards[1278]}), .top({trees[1279], lumberyards[1279]}), .top_right({trees[1280], lumberyards[1280]}), .left({trees[1328], lumberyards[1328]}), .right({trees[1330], lumberyards[1330]}), .bottom_left({trees[1378], lumberyards[1378]}), .bottom({trees[1379], lumberyards[1379]}), .bottom_right({trees[1380], lumberyards[1380]}), .init(2'b00), .state({trees[1329], lumberyards[1329]}));
acre acre_26_30 (.clk(clk), .en(en), .top_left({trees[1279], lumberyards[1279]}), .top({trees[1280], lumberyards[1280]}), .top_right({trees[1281], lumberyards[1281]}), .left({trees[1329], lumberyards[1329]}), .right({trees[1331], lumberyards[1331]}), .bottom_left({trees[1379], lumberyards[1379]}), .bottom({trees[1380], lumberyards[1380]}), .bottom_right({trees[1381], lumberyards[1381]}), .init(2'b00), .state({trees[1330], lumberyards[1330]}));
acre acre_26_31 (.clk(clk), .en(en), .top_left({trees[1280], lumberyards[1280]}), .top({trees[1281], lumberyards[1281]}), .top_right({trees[1282], lumberyards[1282]}), .left({trees[1330], lumberyards[1330]}), .right({trees[1332], lumberyards[1332]}), .bottom_left({trees[1380], lumberyards[1380]}), .bottom({trees[1381], lumberyards[1381]}), .bottom_right({trees[1382], lumberyards[1382]}), .init(2'b00), .state({trees[1331], lumberyards[1331]}));
acre acre_26_32 (.clk(clk), .en(en), .top_left({trees[1281], lumberyards[1281]}), .top({trees[1282], lumberyards[1282]}), .top_right({trees[1283], lumberyards[1283]}), .left({trees[1331], lumberyards[1331]}), .right({trees[1333], lumberyards[1333]}), .bottom_left({trees[1381], lumberyards[1381]}), .bottom({trees[1382], lumberyards[1382]}), .bottom_right({trees[1383], lumberyards[1383]}), .init(2'b00), .state({trees[1332], lumberyards[1332]}));
acre acre_26_33 (.clk(clk), .en(en), .top_left({trees[1282], lumberyards[1282]}), .top({trees[1283], lumberyards[1283]}), .top_right({trees[1284], lumberyards[1284]}), .left({trees[1332], lumberyards[1332]}), .right({trees[1334], lumberyards[1334]}), .bottom_left({trees[1382], lumberyards[1382]}), .bottom({trees[1383], lumberyards[1383]}), .bottom_right({trees[1384], lumberyards[1384]}), .init(2'b00), .state({trees[1333], lumberyards[1333]}));
acre acre_26_34 (.clk(clk), .en(en), .top_left({trees[1283], lumberyards[1283]}), .top({trees[1284], lumberyards[1284]}), .top_right({trees[1285], lumberyards[1285]}), .left({trees[1333], lumberyards[1333]}), .right({trees[1335], lumberyards[1335]}), .bottom_left({trees[1383], lumberyards[1383]}), .bottom({trees[1384], lumberyards[1384]}), .bottom_right({trees[1385], lumberyards[1385]}), .init(2'b10), .state({trees[1334], lumberyards[1334]}));
acre acre_26_35 (.clk(clk), .en(en), .top_left({trees[1284], lumberyards[1284]}), .top({trees[1285], lumberyards[1285]}), .top_right({trees[1286], lumberyards[1286]}), .left({trees[1334], lumberyards[1334]}), .right({trees[1336], lumberyards[1336]}), .bottom_left({trees[1384], lumberyards[1384]}), .bottom({trees[1385], lumberyards[1385]}), .bottom_right({trees[1386], lumberyards[1386]}), .init(2'b01), .state({trees[1335], lumberyards[1335]}));
acre acre_26_36 (.clk(clk), .en(en), .top_left({trees[1285], lumberyards[1285]}), .top({trees[1286], lumberyards[1286]}), .top_right({trees[1287], lumberyards[1287]}), .left({trees[1335], lumberyards[1335]}), .right({trees[1337], lumberyards[1337]}), .bottom_left({trees[1385], lumberyards[1385]}), .bottom({trees[1386], lumberyards[1386]}), .bottom_right({trees[1387], lumberyards[1387]}), .init(2'b00), .state({trees[1336], lumberyards[1336]}));
acre acre_26_37 (.clk(clk), .en(en), .top_left({trees[1286], lumberyards[1286]}), .top({trees[1287], lumberyards[1287]}), .top_right({trees[1288], lumberyards[1288]}), .left({trees[1336], lumberyards[1336]}), .right({trees[1338], lumberyards[1338]}), .bottom_left({trees[1386], lumberyards[1386]}), .bottom({trees[1387], lumberyards[1387]}), .bottom_right({trees[1388], lumberyards[1388]}), .init(2'b00), .state({trees[1337], lumberyards[1337]}));
acre acre_26_38 (.clk(clk), .en(en), .top_left({trees[1287], lumberyards[1287]}), .top({trees[1288], lumberyards[1288]}), .top_right({trees[1289], lumberyards[1289]}), .left({trees[1337], lumberyards[1337]}), .right({trees[1339], lumberyards[1339]}), .bottom_left({trees[1387], lumberyards[1387]}), .bottom({trees[1388], lumberyards[1388]}), .bottom_right({trees[1389], lumberyards[1389]}), .init(2'b10), .state({trees[1338], lumberyards[1338]}));
acre acre_26_39 (.clk(clk), .en(en), .top_left({trees[1288], lumberyards[1288]}), .top({trees[1289], lumberyards[1289]}), .top_right({trees[1290], lumberyards[1290]}), .left({trees[1338], lumberyards[1338]}), .right({trees[1340], lumberyards[1340]}), .bottom_left({trees[1388], lumberyards[1388]}), .bottom({trees[1389], lumberyards[1389]}), .bottom_right({trees[1390], lumberyards[1390]}), .init(2'b00), .state({trees[1339], lumberyards[1339]}));
acre acre_26_40 (.clk(clk), .en(en), .top_left({trees[1289], lumberyards[1289]}), .top({trees[1290], lumberyards[1290]}), .top_right({trees[1291], lumberyards[1291]}), .left({trees[1339], lumberyards[1339]}), .right({trees[1341], lumberyards[1341]}), .bottom_left({trees[1389], lumberyards[1389]}), .bottom({trees[1390], lumberyards[1390]}), .bottom_right({trees[1391], lumberyards[1391]}), .init(2'b01), .state({trees[1340], lumberyards[1340]}));
acre acre_26_41 (.clk(clk), .en(en), .top_left({trees[1290], lumberyards[1290]}), .top({trees[1291], lumberyards[1291]}), .top_right({trees[1292], lumberyards[1292]}), .left({trees[1340], lumberyards[1340]}), .right({trees[1342], lumberyards[1342]}), .bottom_left({trees[1390], lumberyards[1390]}), .bottom({trees[1391], lumberyards[1391]}), .bottom_right({trees[1392], lumberyards[1392]}), .init(2'b00), .state({trees[1341], lumberyards[1341]}));
acre acre_26_42 (.clk(clk), .en(en), .top_left({trees[1291], lumberyards[1291]}), .top({trees[1292], lumberyards[1292]}), .top_right({trees[1293], lumberyards[1293]}), .left({trees[1341], lumberyards[1341]}), .right({trees[1343], lumberyards[1343]}), .bottom_left({trees[1391], lumberyards[1391]}), .bottom({trees[1392], lumberyards[1392]}), .bottom_right({trees[1393], lumberyards[1393]}), .init(2'b00), .state({trees[1342], lumberyards[1342]}));
acre acre_26_43 (.clk(clk), .en(en), .top_left({trees[1292], lumberyards[1292]}), .top({trees[1293], lumberyards[1293]}), .top_right({trees[1294], lumberyards[1294]}), .left({trees[1342], lumberyards[1342]}), .right({trees[1344], lumberyards[1344]}), .bottom_left({trees[1392], lumberyards[1392]}), .bottom({trees[1393], lumberyards[1393]}), .bottom_right({trees[1394], lumberyards[1394]}), .init(2'b00), .state({trees[1343], lumberyards[1343]}));
acre acre_26_44 (.clk(clk), .en(en), .top_left({trees[1293], lumberyards[1293]}), .top({trees[1294], lumberyards[1294]}), .top_right({trees[1295], lumberyards[1295]}), .left({trees[1343], lumberyards[1343]}), .right({trees[1345], lumberyards[1345]}), .bottom_left({trees[1393], lumberyards[1393]}), .bottom({trees[1394], lumberyards[1394]}), .bottom_right({trees[1395], lumberyards[1395]}), .init(2'b00), .state({trees[1344], lumberyards[1344]}));
acre acre_26_45 (.clk(clk), .en(en), .top_left({trees[1294], lumberyards[1294]}), .top({trees[1295], lumberyards[1295]}), .top_right({trees[1296], lumberyards[1296]}), .left({trees[1344], lumberyards[1344]}), .right({trees[1346], lumberyards[1346]}), .bottom_left({trees[1394], lumberyards[1394]}), .bottom({trees[1395], lumberyards[1395]}), .bottom_right({trees[1396], lumberyards[1396]}), .init(2'b01), .state({trees[1345], lumberyards[1345]}));
acre acre_26_46 (.clk(clk), .en(en), .top_left({trees[1295], lumberyards[1295]}), .top({trees[1296], lumberyards[1296]}), .top_right({trees[1297], lumberyards[1297]}), .left({trees[1345], lumberyards[1345]}), .right({trees[1347], lumberyards[1347]}), .bottom_left({trees[1395], lumberyards[1395]}), .bottom({trees[1396], lumberyards[1396]}), .bottom_right({trees[1397], lumberyards[1397]}), .init(2'b00), .state({trees[1346], lumberyards[1346]}));
acre acre_26_47 (.clk(clk), .en(en), .top_left({trees[1296], lumberyards[1296]}), .top({trees[1297], lumberyards[1297]}), .top_right({trees[1298], lumberyards[1298]}), .left({trees[1346], lumberyards[1346]}), .right({trees[1348], lumberyards[1348]}), .bottom_left({trees[1396], lumberyards[1396]}), .bottom({trees[1397], lumberyards[1397]}), .bottom_right({trees[1398], lumberyards[1398]}), .init(2'b00), .state({trees[1347], lumberyards[1347]}));
acre acre_26_48 (.clk(clk), .en(en), .top_left({trees[1297], lumberyards[1297]}), .top({trees[1298], lumberyards[1298]}), .top_right({trees[1299], lumberyards[1299]}), .left({trees[1347], lumberyards[1347]}), .right({trees[1349], lumberyards[1349]}), .bottom_left({trees[1397], lumberyards[1397]}), .bottom({trees[1398], lumberyards[1398]}), .bottom_right({trees[1399], lumberyards[1399]}), .init(2'b01), .state({trees[1348], lumberyards[1348]}));
acre acre_26_49 (.clk(clk), .en(en), .top_left({trees[1298], lumberyards[1298]}), .top({trees[1299], lumberyards[1299]}), .top_right(2'b0), .left({trees[1348], lumberyards[1348]}), .right(2'b0), .bottom_left({trees[1398], lumberyards[1398]}), .bottom({trees[1399], lumberyards[1399]}), .bottom_right(2'b0), .init(2'b00), .state({trees[1349], lumberyards[1349]}));
acre acre_27_0 (.clk(clk), .en(en), .top_left(2'b0), .top({trees[1300], lumberyards[1300]}), .top_right({trees[1301], lumberyards[1301]}), .left(2'b0), .right({trees[1351], lumberyards[1351]}), .bottom_left(2'b0), .bottom({trees[1400], lumberyards[1400]}), .bottom_right({trees[1401], lumberyards[1401]}), .init(2'b10), .state({trees[1350], lumberyards[1350]}));
acre acre_27_1 (.clk(clk), .en(en), .top_left({trees[1300], lumberyards[1300]}), .top({trees[1301], lumberyards[1301]}), .top_right({trees[1302], lumberyards[1302]}), .left({trees[1350], lumberyards[1350]}), .right({trees[1352], lumberyards[1352]}), .bottom_left({trees[1400], lumberyards[1400]}), .bottom({trees[1401], lumberyards[1401]}), .bottom_right({trees[1402], lumberyards[1402]}), .init(2'b01), .state({trees[1351], lumberyards[1351]}));
acre acre_27_2 (.clk(clk), .en(en), .top_left({trees[1301], lumberyards[1301]}), .top({trees[1302], lumberyards[1302]}), .top_right({trees[1303], lumberyards[1303]}), .left({trees[1351], lumberyards[1351]}), .right({trees[1353], lumberyards[1353]}), .bottom_left({trees[1401], lumberyards[1401]}), .bottom({trees[1402], lumberyards[1402]}), .bottom_right({trees[1403], lumberyards[1403]}), .init(2'b00), .state({trees[1352], lumberyards[1352]}));
acre acre_27_3 (.clk(clk), .en(en), .top_left({trees[1302], lumberyards[1302]}), .top({trees[1303], lumberyards[1303]}), .top_right({trees[1304], lumberyards[1304]}), .left({trees[1352], lumberyards[1352]}), .right({trees[1354], lumberyards[1354]}), .bottom_left({trees[1402], lumberyards[1402]}), .bottom({trees[1403], lumberyards[1403]}), .bottom_right({trees[1404], lumberyards[1404]}), .init(2'b00), .state({trees[1353], lumberyards[1353]}));
acre acre_27_4 (.clk(clk), .en(en), .top_left({trees[1303], lumberyards[1303]}), .top({trees[1304], lumberyards[1304]}), .top_right({trees[1305], lumberyards[1305]}), .left({trees[1353], lumberyards[1353]}), .right({trees[1355], lumberyards[1355]}), .bottom_left({trees[1403], lumberyards[1403]}), .bottom({trees[1404], lumberyards[1404]}), .bottom_right({trees[1405], lumberyards[1405]}), .init(2'b01), .state({trees[1354], lumberyards[1354]}));
acre acre_27_5 (.clk(clk), .en(en), .top_left({trees[1304], lumberyards[1304]}), .top({trees[1305], lumberyards[1305]}), .top_right({trees[1306], lumberyards[1306]}), .left({trees[1354], lumberyards[1354]}), .right({trees[1356], lumberyards[1356]}), .bottom_left({trees[1404], lumberyards[1404]}), .bottom({trees[1405], lumberyards[1405]}), .bottom_right({trees[1406], lumberyards[1406]}), .init(2'b00), .state({trees[1355], lumberyards[1355]}));
acre acre_27_6 (.clk(clk), .en(en), .top_left({trees[1305], lumberyards[1305]}), .top({trees[1306], lumberyards[1306]}), .top_right({trees[1307], lumberyards[1307]}), .left({trees[1355], lumberyards[1355]}), .right({trees[1357], lumberyards[1357]}), .bottom_left({trees[1405], lumberyards[1405]}), .bottom({trees[1406], lumberyards[1406]}), .bottom_right({trees[1407], lumberyards[1407]}), .init(2'b00), .state({trees[1356], lumberyards[1356]}));
acre acre_27_7 (.clk(clk), .en(en), .top_left({trees[1306], lumberyards[1306]}), .top({trees[1307], lumberyards[1307]}), .top_right({trees[1308], lumberyards[1308]}), .left({trees[1356], lumberyards[1356]}), .right({trees[1358], lumberyards[1358]}), .bottom_left({trees[1406], lumberyards[1406]}), .bottom({trees[1407], lumberyards[1407]}), .bottom_right({trees[1408], lumberyards[1408]}), .init(2'b01), .state({trees[1357], lumberyards[1357]}));
acre acre_27_8 (.clk(clk), .en(en), .top_left({trees[1307], lumberyards[1307]}), .top({trees[1308], lumberyards[1308]}), .top_right({trees[1309], lumberyards[1309]}), .left({trees[1357], lumberyards[1357]}), .right({trees[1359], lumberyards[1359]}), .bottom_left({trees[1407], lumberyards[1407]}), .bottom({trees[1408], lumberyards[1408]}), .bottom_right({trees[1409], lumberyards[1409]}), .init(2'b01), .state({trees[1358], lumberyards[1358]}));
acre acre_27_9 (.clk(clk), .en(en), .top_left({trees[1308], lumberyards[1308]}), .top({trees[1309], lumberyards[1309]}), .top_right({trees[1310], lumberyards[1310]}), .left({trees[1358], lumberyards[1358]}), .right({trees[1360], lumberyards[1360]}), .bottom_left({trees[1408], lumberyards[1408]}), .bottom({trees[1409], lumberyards[1409]}), .bottom_right({trees[1410], lumberyards[1410]}), .init(2'b00), .state({trees[1359], lumberyards[1359]}));
acre acre_27_10 (.clk(clk), .en(en), .top_left({trees[1309], lumberyards[1309]}), .top({trees[1310], lumberyards[1310]}), .top_right({trees[1311], lumberyards[1311]}), .left({trees[1359], lumberyards[1359]}), .right({trees[1361], lumberyards[1361]}), .bottom_left({trees[1409], lumberyards[1409]}), .bottom({trees[1410], lumberyards[1410]}), .bottom_right({trees[1411], lumberyards[1411]}), .init(2'b00), .state({trees[1360], lumberyards[1360]}));
acre acre_27_11 (.clk(clk), .en(en), .top_left({trees[1310], lumberyards[1310]}), .top({trees[1311], lumberyards[1311]}), .top_right({trees[1312], lumberyards[1312]}), .left({trees[1360], lumberyards[1360]}), .right({trees[1362], lumberyards[1362]}), .bottom_left({trees[1410], lumberyards[1410]}), .bottom({trees[1411], lumberyards[1411]}), .bottom_right({trees[1412], lumberyards[1412]}), .init(2'b00), .state({trees[1361], lumberyards[1361]}));
acre acre_27_12 (.clk(clk), .en(en), .top_left({trees[1311], lumberyards[1311]}), .top({trees[1312], lumberyards[1312]}), .top_right({trees[1313], lumberyards[1313]}), .left({trees[1361], lumberyards[1361]}), .right({trees[1363], lumberyards[1363]}), .bottom_left({trees[1411], lumberyards[1411]}), .bottom({trees[1412], lumberyards[1412]}), .bottom_right({trees[1413], lumberyards[1413]}), .init(2'b00), .state({trees[1362], lumberyards[1362]}));
acre acre_27_13 (.clk(clk), .en(en), .top_left({trees[1312], lumberyards[1312]}), .top({trees[1313], lumberyards[1313]}), .top_right({trees[1314], lumberyards[1314]}), .left({trees[1362], lumberyards[1362]}), .right({trees[1364], lumberyards[1364]}), .bottom_left({trees[1412], lumberyards[1412]}), .bottom({trees[1413], lumberyards[1413]}), .bottom_right({trees[1414], lumberyards[1414]}), .init(2'b00), .state({trees[1363], lumberyards[1363]}));
acre acre_27_14 (.clk(clk), .en(en), .top_left({trees[1313], lumberyards[1313]}), .top({trees[1314], lumberyards[1314]}), .top_right({trees[1315], lumberyards[1315]}), .left({trees[1363], lumberyards[1363]}), .right({trees[1365], lumberyards[1365]}), .bottom_left({trees[1413], lumberyards[1413]}), .bottom({trees[1414], lumberyards[1414]}), .bottom_right({trees[1415], lumberyards[1415]}), .init(2'b01), .state({trees[1364], lumberyards[1364]}));
acre acre_27_15 (.clk(clk), .en(en), .top_left({trees[1314], lumberyards[1314]}), .top({trees[1315], lumberyards[1315]}), .top_right({trees[1316], lumberyards[1316]}), .left({trees[1364], lumberyards[1364]}), .right({trees[1366], lumberyards[1366]}), .bottom_left({trees[1414], lumberyards[1414]}), .bottom({trees[1415], lumberyards[1415]}), .bottom_right({trees[1416], lumberyards[1416]}), .init(2'b10), .state({trees[1365], lumberyards[1365]}));
acre acre_27_16 (.clk(clk), .en(en), .top_left({trees[1315], lumberyards[1315]}), .top({trees[1316], lumberyards[1316]}), .top_right({trees[1317], lumberyards[1317]}), .left({trees[1365], lumberyards[1365]}), .right({trees[1367], lumberyards[1367]}), .bottom_left({trees[1415], lumberyards[1415]}), .bottom({trees[1416], lumberyards[1416]}), .bottom_right({trees[1417], lumberyards[1417]}), .init(2'b01), .state({trees[1366], lumberyards[1366]}));
acre acre_27_17 (.clk(clk), .en(en), .top_left({trees[1316], lumberyards[1316]}), .top({trees[1317], lumberyards[1317]}), .top_right({trees[1318], lumberyards[1318]}), .left({trees[1366], lumberyards[1366]}), .right({trees[1368], lumberyards[1368]}), .bottom_left({trees[1416], lumberyards[1416]}), .bottom({trees[1417], lumberyards[1417]}), .bottom_right({trees[1418], lumberyards[1418]}), .init(2'b10), .state({trees[1367], lumberyards[1367]}));
acre acre_27_18 (.clk(clk), .en(en), .top_left({trees[1317], lumberyards[1317]}), .top({trees[1318], lumberyards[1318]}), .top_right({trees[1319], lumberyards[1319]}), .left({trees[1367], lumberyards[1367]}), .right({trees[1369], lumberyards[1369]}), .bottom_left({trees[1417], lumberyards[1417]}), .bottom({trees[1418], lumberyards[1418]}), .bottom_right({trees[1419], lumberyards[1419]}), .init(2'b00), .state({trees[1368], lumberyards[1368]}));
acre acre_27_19 (.clk(clk), .en(en), .top_left({trees[1318], lumberyards[1318]}), .top({trees[1319], lumberyards[1319]}), .top_right({trees[1320], lumberyards[1320]}), .left({trees[1368], lumberyards[1368]}), .right({trees[1370], lumberyards[1370]}), .bottom_left({trees[1418], lumberyards[1418]}), .bottom({trees[1419], lumberyards[1419]}), .bottom_right({trees[1420], lumberyards[1420]}), .init(2'b00), .state({trees[1369], lumberyards[1369]}));
acre acre_27_20 (.clk(clk), .en(en), .top_left({trees[1319], lumberyards[1319]}), .top({trees[1320], lumberyards[1320]}), .top_right({trees[1321], lumberyards[1321]}), .left({trees[1369], lumberyards[1369]}), .right({trees[1371], lumberyards[1371]}), .bottom_left({trees[1419], lumberyards[1419]}), .bottom({trees[1420], lumberyards[1420]}), .bottom_right({trees[1421], lumberyards[1421]}), .init(2'b00), .state({trees[1370], lumberyards[1370]}));
acre acre_27_21 (.clk(clk), .en(en), .top_left({trees[1320], lumberyards[1320]}), .top({trees[1321], lumberyards[1321]}), .top_right({trees[1322], lumberyards[1322]}), .left({trees[1370], lumberyards[1370]}), .right({trees[1372], lumberyards[1372]}), .bottom_left({trees[1420], lumberyards[1420]}), .bottom({trees[1421], lumberyards[1421]}), .bottom_right({trees[1422], lumberyards[1422]}), .init(2'b01), .state({trees[1371], lumberyards[1371]}));
acre acre_27_22 (.clk(clk), .en(en), .top_left({trees[1321], lumberyards[1321]}), .top({trees[1322], lumberyards[1322]}), .top_right({trees[1323], lumberyards[1323]}), .left({trees[1371], lumberyards[1371]}), .right({trees[1373], lumberyards[1373]}), .bottom_left({trees[1421], lumberyards[1421]}), .bottom({trees[1422], lumberyards[1422]}), .bottom_right({trees[1423], lumberyards[1423]}), .init(2'b00), .state({trees[1372], lumberyards[1372]}));
acre acre_27_23 (.clk(clk), .en(en), .top_left({trees[1322], lumberyards[1322]}), .top({trees[1323], lumberyards[1323]}), .top_right({trees[1324], lumberyards[1324]}), .left({trees[1372], lumberyards[1372]}), .right({trees[1374], lumberyards[1374]}), .bottom_left({trees[1422], lumberyards[1422]}), .bottom({trees[1423], lumberyards[1423]}), .bottom_right({trees[1424], lumberyards[1424]}), .init(2'b00), .state({trees[1373], lumberyards[1373]}));
acre acre_27_24 (.clk(clk), .en(en), .top_left({trees[1323], lumberyards[1323]}), .top({trees[1324], lumberyards[1324]}), .top_right({trees[1325], lumberyards[1325]}), .left({trees[1373], lumberyards[1373]}), .right({trees[1375], lumberyards[1375]}), .bottom_left({trees[1423], lumberyards[1423]}), .bottom({trees[1424], lumberyards[1424]}), .bottom_right({trees[1425], lumberyards[1425]}), .init(2'b00), .state({trees[1374], lumberyards[1374]}));
acre acre_27_25 (.clk(clk), .en(en), .top_left({trees[1324], lumberyards[1324]}), .top({trees[1325], lumberyards[1325]}), .top_right({trees[1326], lumberyards[1326]}), .left({trees[1374], lumberyards[1374]}), .right({trees[1376], lumberyards[1376]}), .bottom_left({trees[1424], lumberyards[1424]}), .bottom({trees[1425], lumberyards[1425]}), .bottom_right({trees[1426], lumberyards[1426]}), .init(2'b00), .state({trees[1375], lumberyards[1375]}));
acre acre_27_26 (.clk(clk), .en(en), .top_left({trees[1325], lumberyards[1325]}), .top({trees[1326], lumberyards[1326]}), .top_right({trees[1327], lumberyards[1327]}), .left({trees[1375], lumberyards[1375]}), .right({trees[1377], lumberyards[1377]}), .bottom_left({trees[1425], lumberyards[1425]}), .bottom({trees[1426], lumberyards[1426]}), .bottom_right({trees[1427], lumberyards[1427]}), .init(2'b00), .state({trees[1376], lumberyards[1376]}));
acre acre_27_27 (.clk(clk), .en(en), .top_left({trees[1326], lumberyards[1326]}), .top({trees[1327], lumberyards[1327]}), .top_right({trees[1328], lumberyards[1328]}), .left({trees[1376], lumberyards[1376]}), .right({trees[1378], lumberyards[1378]}), .bottom_left({trees[1426], lumberyards[1426]}), .bottom({trees[1427], lumberyards[1427]}), .bottom_right({trees[1428], lumberyards[1428]}), .init(2'b01), .state({trees[1377], lumberyards[1377]}));
acre acre_27_28 (.clk(clk), .en(en), .top_left({trees[1327], lumberyards[1327]}), .top({trees[1328], lumberyards[1328]}), .top_right({trees[1329], lumberyards[1329]}), .left({trees[1377], lumberyards[1377]}), .right({trees[1379], lumberyards[1379]}), .bottom_left({trees[1427], lumberyards[1427]}), .bottom({trees[1428], lumberyards[1428]}), .bottom_right({trees[1429], lumberyards[1429]}), .init(2'b00), .state({trees[1378], lumberyards[1378]}));
acre acre_27_29 (.clk(clk), .en(en), .top_left({trees[1328], lumberyards[1328]}), .top({trees[1329], lumberyards[1329]}), .top_right({trees[1330], lumberyards[1330]}), .left({trees[1378], lumberyards[1378]}), .right({trees[1380], lumberyards[1380]}), .bottom_left({trees[1428], lumberyards[1428]}), .bottom({trees[1429], lumberyards[1429]}), .bottom_right({trees[1430], lumberyards[1430]}), .init(2'b00), .state({trees[1379], lumberyards[1379]}));
acre acre_27_30 (.clk(clk), .en(en), .top_left({trees[1329], lumberyards[1329]}), .top({trees[1330], lumberyards[1330]}), .top_right({trees[1331], lumberyards[1331]}), .left({trees[1379], lumberyards[1379]}), .right({trees[1381], lumberyards[1381]}), .bottom_left({trees[1429], lumberyards[1429]}), .bottom({trees[1430], lumberyards[1430]}), .bottom_right({trees[1431], lumberyards[1431]}), .init(2'b00), .state({trees[1380], lumberyards[1380]}));
acre acre_27_31 (.clk(clk), .en(en), .top_left({trees[1330], lumberyards[1330]}), .top({trees[1331], lumberyards[1331]}), .top_right({trees[1332], lumberyards[1332]}), .left({trees[1380], lumberyards[1380]}), .right({trees[1382], lumberyards[1382]}), .bottom_left({trees[1430], lumberyards[1430]}), .bottom({trees[1431], lumberyards[1431]}), .bottom_right({trees[1432], lumberyards[1432]}), .init(2'b00), .state({trees[1381], lumberyards[1381]}));
acre acre_27_32 (.clk(clk), .en(en), .top_left({trees[1331], lumberyards[1331]}), .top({trees[1332], lumberyards[1332]}), .top_right({trees[1333], lumberyards[1333]}), .left({trees[1381], lumberyards[1381]}), .right({trees[1383], lumberyards[1383]}), .bottom_left({trees[1431], lumberyards[1431]}), .bottom({trees[1432], lumberyards[1432]}), .bottom_right({trees[1433], lumberyards[1433]}), .init(2'b10), .state({trees[1382], lumberyards[1382]}));
acre acre_27_33 (.clk(clk), .en(en), .top_left({trees[1332], lumberyards[1332]}), .top({trees[1333], lumberyards[1333]}), .top_right({trees[1334], lumberyards[1334]}), .left({trees[1382], lumberyards[1382]}), .right({trees[1384], lumberyards[1384]}), .bottom_left({trees[1432], lumberyards[1432]}), .bottom({trees[1433], lumberyards[1433]}), .bottom_right({trees[1434], lumberyards[1434]}), .init(2'b00), .state({trees[1383], lumberyards[1383]}));
acre acre_27_34 (.clk(clk), .en(en), .top_left({trees[1333], lumberyards[1333]}), .top({trees[1334], lumberyards[1334]}), .top_right({trees[1335], lumberyards[1335]}), .left({trees[1383], lumberyards[1383]}), .right({trees[1385], lumberyards[1385]}), .bottom_left({trees[1433], lumberyards[1433]}), .bottom({trees[1434], lumberyards[1434]}), .bottom_right({trees[1435], lumberyards[1435]}), .init(2'b10), .state({trees[1384], lumberyards[1384]}));
acre acre_27_35 (.clk(clk), .en(en), .top_left({trees[1334], lumberyards[1334]}), .top({trees[1335], lumberyards[1335]}), .top_right({trees[1336], lumberyards[1336]}), .left({trees[1384], lumberyards[1384]}), .right({trees[1386], lumberyards[1386]}), .bottom_left({trees[1434], lumberyards[1434]}), .bottom({trees[1435], lumberyards[1435]}), .bottom_right({trees[1436], lumberyards[1436]}), .init(2'b00), .state({trees[1385], lumberyards[1385]}));
acre acre_27_36 (.clk(clk), .en(en), .top_left({trees[1335], lumberyards[1335]}), .top({trees[1336], lumberyards[1336]}), .top_right({trees[1337], lumberyards[1337]}), .left({trees[1385], lumberyards[1385]}), .right({trees[1387], lumberyards[1387]}), .bottom_left({trees[1435], lumberyards[1435]}), .bottom({trees[1436], lumberyards[1436]}), .bottom_right({trees[1437], lumberyards[1437]}), .init(2'b10), .state({trees[1386], lumberyards[1386]}));
acre acre_27_37 (.clk(clk), .en(en), .top_left({trees[1336], lumberyards[1336]}), .top({trees[1337], lumberyards[1337]}), .top_right({trees[1338], lumberyards[1338]}), .left({trees[1386], lumberyards[1386]}), .right({trees[1388], lumberyards[1388]}), .bottom_left({trees[1436], lumberyards[1436]}), .bottom({trees[1437], lumberyards[1437]}), .bottom_right({trees[1438], lumberyards[1438]}), .init(2'b00), .state({trees[1387], lumberyards[1387]}));
acre acre_27_38 (.clk(clk), .en(en), .top_left({trees[1337], lumberyards[1337]}), .top({trees[1338], lumberyards[1338]}), .top_right({trees[1339], lumberyards[1339]}), .left({trees[1387], lumberyards[1387]}), .right({trees[1389], lumberyards[1389]}), .bottom_left({trees[1437], lumberyards[1437]}), .bottom({trees[1438], lumberyards[1438]}), .bottom_right({trees[1439], lumberyards[1439]}), .init(2'b00), .state({trees[1388], lumberyards[1388]}));
acre acre_27_39 (.clk(clk), .en(en), .top_left({trees[1338], lumberyards[1338]}), .top({trees[1339], lumberyards[1339]}), .top_right({trees[1340], lumberyards[1340]}), .left({trees[1388], lumberyards[1388]}), .right({trees[1390], lumberyards[1390]}), .bottom_left({trees[1438], lumberyards[1438]}), .bottom({trees[1439], lumberyards[1439]}), .bottom_right({trees[1440], lumberyards[1440]}), .init(2'b10), .state({trees[1389], lumberyards[1389]}));
acre acre_27_40 (.clk(clk), .en(en), .top_left({trees[1339], lumberyards[1339]}), .top({trees[1340], lumberyards[1340]}), .top_right({trees[1341], lumberyards[1341]}), .left({trees[1389], lumberyards[1389]}), .right({trees[1391], lumberyards[1391]}), .bottom_left({trees[1439], lumberyards[1439]}), .bottom({trees[1440], lumberyards[1440]}), .bottom_right({trees[1441], lumberyards[1441]}), .init(2'b00), .state({trees[1390], lumberyards[1390]}));
acre acre_27_41 (.clk(clk), .en(en), .top_left({trees[1340], lumberyards[1340]}), .top({trees[1341], lumberyards[1341]}), .top_right({trees[1342], lumberyards[1342]}), .left({trees[1390], lumberyards[1390]}), .right({trees[1392], lumberyards[1392]}), .bottom_left({trees[1440], lumberyards[1440]}), .bottom({trees[1441], lumberyards[1441]}), .bottom_right({trees[1442], lumberyards[1442]}), .init(2'b00), .state({trees[1391], lumberyards[1391]}));
acre acre_27_42 (.clk(clk), .en(en), .top_left({trees[1341], lumberyards[1341]}), .top({trees[1342], lumberyards[1342]}), .top_right({trees[1343], lumberyards[1343]}), .left({trees[1391], lumberyards[1391]}), .right({trees[1393], lumberyards[1393]}), .bottom_left({trees[1441], lumberyards[1441]}), .bottom({trees[1442], lumberyards[1442]}), .bottom_right({trees[1443], lumberyards[1443]}), .init(2'b01), .state({trees[1392], lumberyards[1392]}));
acre acre_27_43 (.clk(clk), .en(en), .top_left({trees[1342], lumberyards[1342]}), .top({trees[1343], lumberyards[1343]}), .top_right({trees[1344], lumberyards[1344]}), .left({trees[1392], lumberyards[1392]}), .right({trees[1394], lumberyards[1394]}), .bottom_left({trees[1442], lumberyards[1442]}), .bottom({trees[1443], lumberyards[1443]}), .bottom_right({trees[1444], lumberyards[1444]}), .init(2'b00), .state({trees[1393], lumberyards[1393]}));
acre acre_27_44 (.clk(clk), .en(en), .top_left({trees[1343], lumberyards[1343]}), .top({trees[1344], lumberyards[1344]}), .top_right({trees[1345], lumberyards[1345]}), .left({trees[1393], lumberyards[1393]}), .right({trees[1395], lumberyards[1395]}), .bottom_left({trees[1443], lumberyards[1443]}), .bottom({trees[1444], lumberyards[1444]}), .bottom_right({trees[1445], lumberyards[1445]}), .init(2'b10), .state({trees[1394], lumberyards[1394]}));
acre acre_27_45 (.clk(clk), .en(en), .top_left({trees[1344], lumberyards[1344]}), .top({trees[1345], lumberyards[1345]}), .top_right({trees[1346], lumberyards[1346]}), .left({trees[1394], lumberyards[1394]}), .right({trees[1396], lumberyards[1396]}), .bottom_left({trees[1444], lumberyards[1444]}), .bottom({trees[1445], lumberyards[1445]}), .bottom_right({trees[1446], lumberyards[1446]}), .init(2'b00), .state({trees[1395], lumberyards[1395]}));
acre acre_27_46 (.clk(clk), .en(en), .top_left({trees[1345], lumberyards[1345]}), .top({trees[1346], lumberyards[1346]}), .top_right({trees[1347], lumberyards[1347]}), .left({trees[1395], lumberyards[1395]}), .right({trees[1397], lumberyards[1397]}), .bottom_left({trees[1445], lumberyards[1445]}), .bottom({trees[1446], lumberyards[1446]}), .bottom_right({trees[1447], lumberyards[1447]}), .init(2'b00), .state({trees[1396], lumberyards[1396]}));
acre acre_27_47 (.clk(clk), .en(en), .top_left({trees[1346], lumberyards[1346]}), .top({trees[1347], lumberyards[1347]}), .top_right({trees[1348], lumberyards[1348]}), .left({trees[1396], lumberyards[1396]}), .right({trees[1398], lumberyards[1398]}), .bottom_left({trees[1446], lumberyards[1446]}), .bottom({trees[1447], lumberyards[1447]}), .bottom_right({trees[1448], lumberyards[1448]}), .init(2'b01), .state({trees[1397], lumberyards[1397]}));
acre acre_27_48 (.clk(clk), .en(en), .top_left({trees[1347], lumberyards[1347]}), .top({trees[1348], lumberyards[1348]}), .top_right({trees[1349], lumberyards[1349]}), .left({trees[1397], lumberyards[1397]}), .right({trees[1399], lumberyards[1399]}), .bottom_left({trees[1447], lumberyards[1447]}), .bottom({trees[1448], lumberyards[1448]}), .bottom_right({trees[1449], lumberyards[1449]}), .init(2'b10), .state({trees[1398], lumberyards[1398]}));
acre acre_27_49 (.clk(clk), .en(en), .top_left({trees[1348], lumberyards[1348]}), .top({trees[1349], lumberyards[1349]}), .top_right(2'b0), .left({trees[1398], lumberyards[1398]}), .right(2'b0), .bottom_left({trees[1448], lumberyards[1448]}), .bottom({trees[1449], lumberyards[1449]}), .bottom_right(2'b0), .init(2'b00), .state({trees[1399], lumberyards[1399]}));
acre acre_28_0 (.clk(clk), .en(en), .top_left(2'b0), .top({trees[1350], lumberyards[1350]}), .top_right({trees[1351], lumberyards[1351]}), .left(2'b0), .right({trees[1401], lumberyards[1401]}), .bottom_left(2'b0), .bottom({trees[1450], lumberyards[1450]}), .bottom_right({trees[1451], lumberyards[1451]}), .init(2'b00), .state({trees[1400], lumberyards[1400]}));
acre acre_28_1 (.clk(clk), .en(en), .top_left({trees[1350], lumberyards[1350]}), .top({trees[1351], lumberyards[1351]}), .top_right({trees[1352], lumberyards[1352]}), .left({trees[1400], lumberyards[1400]}), .right({trees[1402], lumberyards[1402]}), .bottom_left({trees[1450], lumberyards[1450]}), .bottom({trees[1451], lumberyards[1451]}), .bottom_right({trees[1452], lumberyards[1452]}), .init(2'b01), .state({trees[1401], lumberyards[1401]}));
acre acre_28_2 (.clk(clk), .en(en), .top_left({trees[1351], lumberyards[1351]}), .top({trees[1352], lumberyards[1352]}), .top_right({trees[1353], lumberyards[1353]}), .left({trees[1401], lumberyards[1401]}), .right({trees[1403], lumberyards[1403]}), .bottom_left({trees[1451], lumberyards[1451]}), .bottom({trees[1452], lumberyards[1452]}), .bottom_right({trees[1453], lumberyards[1453]}), .init(2'b00), .state({trees[1402], lumberyards[1402]}));
acre acre_28_3 (.clk(clk), .en(en), .top_left({trees[1352], lumberyards[1352]}), .top({trees[1353], lumberyards[1353]}), .top_right({trees[1354], lumberyards[1354]}), .left({trees[1402], lumberyards[1402]}), .right({trees[1404], lumberyards[1404]}), .bottom_left({trees[1452], lumberyards[1452]}), .bottom({trees[1453], lumberyards[1453]}), .bottom_right({trees[1454], lumberyards[1454]}), .init(2'b01), .state({trees[1403], lumberyards[1403]}));
acre acre_28_4 (.clk(clk), .en(en), .top_left({trees[1353], lumberyards[1353]}), .top({trees[1354], lumberyards[1354]}), .top_right({trees[1355], lumberyards[1355]}), .left({trees[1403], lumberyards[1403]}), .right({trees[1405], lumberyards[1405]}), .bottom_left({trees[1453], lumberyards[1453]}), .bottom({trees[1454], lumberyards[1454]}), .bottom_right({trees[1455], lumberyards[1455]}), .init(2'b10), .state({trees[1404], lumberyards[1404]}));
acre acre_28_5 (.clk(clk), .en(en), .top_left({trees[1354], lumberyards[1354]}), .top({trees[1355], lumberyards[1355]}), .top_right({trees[1356], lumberyards[1356]}), .left({trees[1404], lumberyards[1404]}), .right({trees[1406], lumberyards[1406]}), .bottom_left({trees[1454], lumberyards[1454]}), .bottom({trees[1455], lumberyards[1455]}), .bottom_right({trees[1456], lumberyards[1456]}), .init(2'b01), .state({trees[1405], lumberyards[1405]}));
acre acre_28_6 (.clk(clk), .en(en), .top_left({trees[1355], lumberyards[1355]}), .top({trees[1356], lumberyards[1356]}), .top_right({trees[1357], lumberyards[1357]}), .left({trees[1405], lumberyards[1405]}), .right({trees[1407], lumberyards[1407]}), .bottom_left({trees[1455], lumberyards[1455]}), .bottom({trees[1456], lumberyards[1456]}), .bottom_right({trees[1457], lumberyards[1457]}), .init(2'b00), .state({trees[1406], lumberyards[1406]}));
acre acre_28_7 (.clk(clk), .en(en), .top_left({trees[1356], lumberyards[1356]}), .top({trees[1357], lumberyards[1357]}), .top_right({trees[1358], lumberyards[1358]}), .left({trees[1406], lumberyards[1406]}), .right({trees[1408], lumberyards[1408]}), .bottom_left({trees[1456], lumberyards[1456]}), .bottom({trees[1457], lumberyards[1457]}), .bottom_right({trees[1458], lumberyards[1458]}), .init(2'b00), .state({trees[1407], lumberyards[1407]}));
acre acre_28_8 (.clk(clk), .en(en), .top_left({trees[1357], lumberyards[1357]}), .top({trees[1358], lumberyards[1358]}), .top_right({trees[1359], lumberyards[1359]}), .left({trees[1407], lumberyards[1407]}), .right({trees[1409], lumberyards[1409]}), .bottom_left({trees[1457], lumberyards[1457]}), .bottom({trees[1458], lumberyards[1458]}), .bottom_right({trees[1459], lumberyards[1459]}), .init(2'b01), .state({trees[1408], lumberyards[1408]}));
acre acre_28_9 (.clk(clk), .en(en), .top_left({trees[1358], lumberyards[1358]}), .top({trees[1359], lumberyards[1359]}), .top_right({trees[1360], lumberyards[1360]}), .left({trees[1408], lumberyards[1408]}), .right({trees[1410], lumberyards[1410]}), .bottom_left({trees[1458], lumberyards[1458]}), .bottom({trees[1459], lumberyards[1459]}), .bottom_right({trees[1460], lumberyards[1460]}), .init(2'b10), .state({trees[1409], lumberyards[1409]}));
acre acre_28_10 (.clk(clk), .en(en), .top_left({trees[1359], lumberyards[1359]}), .top({trees[1360], lumberyards[1360]}), .top_right({trees[1361], lumberyards[1361]}), .left({trees[1409], lumberyards[1409]}), .right({trees[1411], lumberyards[1411]}), .bottom_left({trees[1459], lumberyards[1459]}), .bottom({trees[1460], lumberyards[1460]}), .bottom_right({trees[1461], lumberyards[1461]}), .init(2'b00), .state({trees[1410], lumberyards[1410]}));
acre acre_28_11 (.clk(clk), .en(en), .top_left({trees[1360], lumberyards[1360]}), .top({trees[1361], lumberyards[1361]}), .top_right({trees[1362], lumberyards[1362]}), .left({trees[1410], lumberyards[1410]}), .right({trees[1412], lumberyards[1412]}), .bottom_left({trees[1460], lumberyards[1460]}), .bottom({trees[1461], lumberyards[1461]}), .bottom_right({trees[1462], lumberyards[1462]}), .init(2'b00), .state({trees[1411], lumberyards[1411]}));
acre acre_28_12 (.clk(clk), .en(en), .top_left({trees[1361], lumberyards[1361]}), .top({trees[1362], lumberyards[1362]}), .top_right({trees[1363], lumberyards[1363]}), .left({trees[1411], lumberyards[1411]}), .right({trees[1413], lumberyards[1413]}), .bottom_left({trees[1461], lumberyards[1461]}), .bottom({trees[1462], lumberyards[1462]}), .bottom_right({trees[1463], lumberyards[1463]}), .init(2'b10), .state({trees[1412], lumberyards[1412]}));
acre acre_28_13 (.clk(clk), .en(en), .top_left({trees[1362], lumberyards[1362]}), .top({trees[1363], lumberyards[1363]}), .top_right({trees[1364], lumberyards[1364]}), .left({trees[1412], lumberyards[1412]}), .right({trees[1414], lumberyards[1414]}), .bottom_left({trees[1462], lumberyards[1462]}), .bottom({trees[1463], lumberyards[1463]}), .bottom_right({trees[1464], lumberyards[1464]}), .init(2'b00), .state({trees[1413], lumberyards[1413]}));
acre acre_28_14 (.clk(clk), .en(en), .top_left({trees[1363], lumberyards[1363]}), .top({trees[1364], lumberyards[1364]}), .top_right({trees[1365], lumberyards[1365]}), .left({trees[1413], lumberyards[1413]}), .right({trees[1415], lumberyards[1415]}), .bottom_left({trees[1463], lumberyards[1463]}), .bottom({trees[1464], lumberyards[1464]}), .bottom_right({trees[1465], lumberyards[1465]}), .init(2'b01), .state({trees[1414], lumberyards[1414]}));
acre acre_28_15 (.clk(clk), .en(en), .top_left({trees[1364], lumberyards[1364]}), .top({trees[1365], lumberyards[1365]}), .top_right({trees[1366], lumberyards[1366]}), .left({trees[1414], lumberyards[1414]}), .right({trees[1416], lumberyards[1416]}), .bottom_left({trees[1464], lumberyards[1464]}), .bottom({trees[1465], lumberyards[1465]}), .bottom_right({trees[1466], lumberyards[1466]}), .init(2'b00), .state({trees[1415], lumberyards[1415]}));
acre acre_28_16 (.clk(clk), .en(en), .top_left({trees[1365], lumberyards[1365]}), .top({trees[1366], lumberyards[1366]}), .top_right({trees[1367], lumberyards[1367]}), .left({trees[1415], lumberyards[1415]}), .right({trees[1417], lumberyards[1417]}), .bottom_left({trees[1465], lumberyards[1465]}), .bottom({trees[1466], lumberyards[1466]}), .bottom_right({trees[1467], lumberyards[1467]}), .init(2'b00), .state({trees[1416], lumberyards[1416]}));
acre acre_28_17 (.clk(clk), .en(en), .top_left({trees[1366], lumberyards[1366]}), .top({trees[1367], lumberyards[1367]}), .top_right({trees[1368], lumberyards[1368]}), .left({trees[1416], lumberyards[1416]}), .right({trees[1418], lumberyards[1418]}), .bottom_left({trees[1466], lumberyards[1466]}), .bottom({trees[1467], lumberyards[1467]}), .bottom_right({trees[1468], lumberyards[1468]}), .init(2'b10), .state({trees[1417], lumberyards[1417]}));
acre acre_28_18 (.clk(clk), .en(en), .top_left({trees[1367], lumberyards[1367]}), .top({trees[1368], lumberyards[1368]}), .top_right({trees[1369], lumberyards[1369]}), .left({trees[1417], lumberyards[1417]}), .right({trees[1419], lumberyards[1419]}), .bottom_left({trees[1467], lumberyards[1467]}), .bottom({trees[1468], lumberyards[1468]}), .bottom_right({trees[1469], lumberyards[1469]}), .init(2'b00), .state({trees[1418], lumberyards[1418]}));
acre acre_28_19 (.clk(clk), .en(en), .top_left({trees[1368], lumberyards[1368]}), .top({trees[1369], lumberyards[1369]}), .top_right({trees[1370], lumberyards[1370]}), .left({trees[1418], lumberyards[1418]}), .right({trees[1420], lumberyards[1420]}), .bottom_left({trees[1468], lumberyards[1468]}), .bottom({trees[1469], lumberyards[1469]}), .bottom_right({trees[1470], lumberyards[1470]}), .init(2'b00), .state({trees[1419], lumberyards[1419]}));
acre acre_28_20 (.clk(clk), .en(en), .top_left({trees[1369], lumberyards[1369]}), .top({trees[1370], lumberyards[1370]}), .top_right({trees[1371], lumberyards[1371]}), .left({trees[1419], lumberyards[1419]}), .right({trees[1421], lumberyards[1421]}), .bottom_left({trees[1469], lumberyards[1469]}), .bottom({trees[1470], lumberyards[1470]}), .bottom_right({trees[1471], lumberyards[1471]}), .init(2'b10), .state({trees[1420], lumberyards[1420]}));
acre acre_28_21 (.clk(clk), .en(en), .top_left({trees[1370], lumberyards[1370]}), .top({trees[1371], lumberyards[1371]}), .top_right({trees[1372], lumberyards[1372]}), .left({trees[1420], lumberyards[1420]}), .right({trees[1422], lumberyards[1422]}), .bottom_left({trees[1470], lumberyards[1470]}), .bottom({trees[1471], lumberyards[1471]}), .bottom_right({trees[1472], lumberyards[1472]}), .init(2'b01), .state({trees[1421], lumberyards[1421]}));
acre acre_28_22 (.clk(clk), .en(en), .top_left({trees[1371], lumberyards[1371]}), .top({trees[1372], lumberyards[1372]}), .top_right({trees[1373], lumberyards[1373]}), .left({trees[1421], lumberyards[1421]}), .right({trees[1423], lumberyards[1423]}), .bottom_left({trees[1471], lumberyards[1471]}), .bottom({trees[1472], lumberyards[1472]}), .bottom_right({trees[1473], lumberyards[1473]}), .init(2'b10), .state({trees[1422], lumberyards[1422]}));
acre acre_28_23 (.clk(clk), .en(en), .top_left({trees[1372], lumberyards[1372]}), .top({trees[1373], lumberyards[1373]}), .top_right({trees[1374], lumberyards[1374]}), .left({trees[1422], lumberyards[1422]}), .right({trees[1424], lumberyards[1424]}), .bottom_left({trees[1472], lumberyards[1472]}), .bottom({trees[1473], lumberyards[1473]}), .bottom_right({trees[1474], lumberyards[1474]}), .init(2'b10), .state({trees[1423], lumberyards[1423]}));
acre acre_28_24 (.clk(clk), .en(en), .top_left({trees[1373], lumberyards[1373]}), .top({trees[1374], lumberyards[1374]}), .top_right({trees[1375], lumberyards[1375]}), .left({trees[1423], lumberyards[1423]}), .right({trees[1425], lumberyards[1425]}), .bottom_left({trees[1473], lumberyards[1473]}), .bottom({trees[1474], lumberyards[1474]}), .bottom_right({trees[1475], lumberyards[1475]}), .init(2'b10), .state({trees[1424], lumberyards[1424]}));
acre acre_28_25 (.clk(clk), .en(en), .top_left({trees[1374], lumberyards[1374]}), .top({trees[1375], lumberyards[1375]}), .top_right({trees[1376], lumberyards[1376]}), .left({trees[1424], lumberyards[1424]}), .right({trees[1426], lumberyards[1426]}), .bottom_left({trees[1474], lumberyards[1474]}), .bottom({trees[1475], lumberyards[1475]}), .bottom_right({trees[1476], lumberyards[1476]}), .init(2'b10), .state({trees[1425], lumberyards[1425]}));
acre acre_28_26 (.clk(clk), .en(en), .top_left({trees[1375], lumberyards[1375]}), .top({trees[1376], lumberyards[1376]}), .top_right({trees[1377], lumberyards[1377]}), .left({trees[1425], lumberyards[1425]}), .right({trees[1427], lumberyards[1427]}), .bottom_left({trees[1475], lumberyards[1475]}), .bottom({trees[1476], lumberyards[1476]}), .bottom_right({trees[1477], lumberyards[1477]}), .init(2'b00), .state({trees[1426], lumberyards[1426]}));
acre acre_28_27 (.clk(clk), .en(en), .top_left({trees[1376], lumberyards[1376]}), .top({trees[1377], lumberyards[1377]}), .top_right({trees[1378], lumberyards[1378]}), .left({trees[1426], lumberyards[1426]}), .right({trees[1428], lumberyards[1428]}), .bottom_left({trees[1476], lumberyards[1476]}), .bottom({trees[1477], lumberyards[1477]}), .bottom_right({trees[1478], lumberyards[1478]}), .init(2'b00), .state({trees[1427], lumberyards[1427]}));
acre acre_28_28 (.clk(clk), .en(en), .top_left({trees[1377], lumberyards[1377]}), .top({trees[1378], lumberyards[1378]}), .top_right({trees[1379], lumberyards[1379]}), .left({trees[1427], lumberyards[1427]}), .right({trees[1429], lumberyards[1429]}), .bottom_left({trees[1477], lumberyards[1477]}), .bottom({trees[1478], lumberyards[1478]}), .bottom_right({trees[1479], lumberyards[1479]}), .init(2'b01), .state({trees[1428], lumberyards[1428]}));
acre acre_28_29 (.clk(clk), .en(en), .top_left({trees[1378], lumberyards[1378]}), .top({trees[1379], lumberyards[1379]}), .top_right({trees[1380], lumberyards[1380]}), .left({trees[1428], lumberyards[1428]}), .right({trees[1430], lumberyards[1430]}), .bottom_left({trees[1478], lumberyards[1478]}), .bottom({trees[1479], lumberyards[1479]}), .bottom_right({trees[1480], lumberyards[1480]}), .init(2'b01), .state({trees[1429], lumberyards[1429]}));
acre acre_28_30 (.clk(clk), .en(en), .top_left({trees[1379], lumberyards[1379]}), .top({trees[1380], lumberyards[1380]}), .top_right({trees[1381], lumberyards[1381]}), .left({trees[1429], lumberyards[1429]}), .right({trees[1431], lumberyards[1431]}), .bottom_left({trees[1479], lumberyards[1479]}), .bottom({trees[1480], lumberyards[1480]}), .bottom_right({trees[1481], lumberyards[1481]}), .init(2'b00), .state({trees[1430], lumberyards[1430]}));
acre acre_28_31 (.clk(clk), .en(en), .top_left({trees[1380], lumberyards[1380]}), .top({trees[1381], lumberyards[1381]}), .top_right({trees[1382], lumberyards[1382]}), .left({trees[1430], lumberyards[1430]}), .right({trees[1432], lumberyards[1432]}), .bottom_left({trees[1480], lumberyards[1480]}), .bottom({trees[1481], lumberyards[1481]}), .bottom_right({trees[1482], lumberyards[1482]}), .init(2'b01), .state({trees[1431], lumberyards[1431]}));
acre acre_28_32 (.clk(clk), .en(en), .top_left({trees[1381], lumberyards[1381]}), .top({trees[1382], lumberyards[1382]}), .top_right({trees[1383], lumberyards[1383]}), .left({trees[1431], lumberyards[1431]}), .right({trees[1433], lumberyards[1433]}), .bottom_left({trees[1481], lumberyards[1481]}), .bottom({trees[1482], lumberyards[1482]}), .bottom_right({trees[1483], lumberyards[1483]}), .init(2'b10), .state({trees[1432], lumberyards[1432]}));
acre acre_28_33 (.clk(clk), .en(en), .top_left({trees[1382], lumberyards[1382]}), .top({trees[1383], lumberyards[1383]}), .top_right({trees[1384], lumberyards[1384]}), .left({trees[1432], lumberyards[1432]}), .right({trees[1434], lumberyards[1434]}), .bottom_left({trees[1482], lumberyards[1482]}), .bottom({trees[1483], lumberyards[1483]}), .bottom_right({trees[1484], lumberyards[1484]}), .init(2'b00), .state({trees[1433], lumberyards[1433]}));
acre acre_28_34 (.clk(clk), .en(en), .top_left({trees[1383], lumberyards[1383]}), .top({trees[1384], lumberyards[1384]}), .top_right({trees[1385], lumberyards[1385]}), .left({trees[1433], lumberyards[1433]}), .right({trees[1435], lumberyards[1435]}), .bottom_left({trees[1483], lumberyards[1483]}), .bottom({trees[1484], lumberyards[1484]}), .bottom_right({trees[1485], lumberyards[1485]}), .init(2'b00), .state({trees[1434], lumberyards[1434]}));
acre acre_28_35 (.clk(clk), .en(en), .top_left({trees[1384], lumberyards[1384]}), .top({trees[1385], lumberyards[1385]}), .top_right({trees[1386], lumberyards[1386]}), .left({trees[1434], lumberyards[1434]}), .right({trees[1436], lumberyards[1436]}), .bottom_left({trees[1484], lumberyards[1484]}), .bottom({trees[1485], lumberyards[1485]}), .bottom_right({trees[1486], lumberyards[1486]}), .init(2'b10), .state({trees[1435], lumberyards[1435]}));
acre acre_28_36 (.clk(clk), .en(en), .top_left({trees[1385], lumberyards[1385]}), .top({trees[1386], lumberyards[1386]}), .top_right({trees[1387], lumberyards[1387]}), .left({trees[1435], lumberyards[1435]}), .right({trees[1437], lumberyards[1437]}), .bottom_left({trees[1485], lumberyards[1485]}), .bottom({trees[1486], lumberyards[1486]}), .bottom_right({trees[1487], lumberyards[1487]}), .init(2'b00), .state({trees[1436], lumberyards[1436]}));
acre acre_28_37 (.clk(clk), .en(en), .top_left({trees[1386], lumberyards[1386]}), .top({trees[1387], lumberyards[1387]}), .top_right({trees[1388], lumberyards[1388]}), .left({trees[1436], lumberyards[1436]}), .right({trees[1438], lumberyards[1438]}), .bottom_left({trees[1486], lumberyards[1486]}), .bottom({trees[1487], lumberyards[1487]}), .bottom_right({trees[1488], lumberyards[1488]}), .init(2'b00), .state({trees[1437], lumberyards[1437]}));
acre acre_28_38 (.clk(clk), .en(en), .top_left({trees[1387], lumberyards[1387]}), .top({trees[1388], lumberyards[1388]}), .top_right({trees[1389], lumberyards[1389]}), .left({trees[1437], lumberyards[1437]}), .right({trees[1439], lumberyards[1439]}), .bottom_left({trees[1487], lumberyards[1487]}), .bottom({trees[1488], lumberyards[1488]}), .bottom_right({trees[1489], lumberyards[1489]}), .init(2'b01), .state({trees[1438], lumberyards[1438]}));
acre acre_28_39 (.clk(clk), .en(en), .top_left({trees[1388], lumberyards[1388]}), .top({trees[1389], lumberyards[1389]}), .top_right({trees[1390], lumberyards[1390]}), .left({trees[1438], lumberyards[1438]}), .right({trees[1440], lumberyards[1440]}), .bottom_left({trees[1488], lumberyards[1488]}), .bottom({trees[1489], lumberyards[1489]}), .bottom_right({trees[1490], lumberyards[1490]}), .init(2'b00), .state({trees[1439], lumberyards[1439]}));
acre acre_28_40 (.clk(clk), .en(en), .top_left({trees[1389], lumberyards[1389]}), .top({trees[1390], lumberyards[1390]}), .top_right({trees[1391], lumberyards[1391]}), .left({trees[1439], lumberyards[1439]}), .right({trees[1441], lumberyards[1441]}), .bottom_left({trees[1489], lumberyards[1489]}), .bottom({trees[1490], lumberyards[1490]}), .bottom_right({trees[1491], lumberyards[1491]}), .init(2'b10), .state({trees[1440], lumberyards[1440]}));
acre acre_28_41 (.clk(clk), .en(en), .top_left({trees[1390], lumberyards[1390]}), .top({trees[1391], lumberyards[1391]}), .top_right({trees[1392], lumberyards[1392]}), .left({trees[1440], lumberyards[1440]}), .right({trees[1442], lumberyards[1442]}), .bottom_left({trees[1490], lumberyards[1490]}), .bottom({trees[1491], lumberyards[1491]}), .bottom_right({trees[1492], lumberyards[1492]}), .init(2'b01), .state({trees[1441], lumberyards[1441]}));
acre acre_28_42 (.clk(clk), .en(en), .top_left({trees[1391], lumberyards[1391]}), .top({trees[1392], lumberyards[1392]}), .top_right({trees[1393], lumberyards[1393]}), .left({trees[1441], lumberyards[1441]}), .right({trees[1443], lumberyards[1443]}), .bottom_left({trees[1491], lumberyards[1491]}), .bottom({trees[1492], lumberyards[1492]}), .bottom_right({trees[1493], lumberyards[1493]}), .init(2'b01), .state({trees[1442], lumberyards[1442]}));
acre acre_28_43 (.clk(clk), .en(en), .top_left({trees[1392], lumberyards[1392]}), .top({trees[1393], lumberyards[1393]}), .top_right({trees[1394], lumberyards[1394]}), .left({trees[1442], lumberyards[1442]}), .right({trees[1444], lumberyards[1444]}), .bottom_left({trees[1492], lumberyards[1492]}), .bottom({trees[1493], lumberyards[1493]}), .bottom_right({trees[1494], lumberyards[1494]}), .init(2'b00), .state({trees[1443], lumberyards[1443]}));
acre acre_28_44 (.clk(clk), .en(en), .top_left({trees[1393], lumberyards[1393]}), .top({trees[1394], lumberyards[1394]}), .top_right({trees[1395], lumberyards[1395]}), .left({trees[1443], lumberyards[1443]}), .right({trees[1445], lumberyards[1445]}), .bottom_left({trees[1493], lumberyards[1493]}), .bottom({trees[1494], lumberyards[1494]}), .bottom_right({trees[1495], lumberyards[1495]}), .init(2'b10), .state({trees[1444], lumberyards[1444]}));
acre acre_28_45 (.clk(clk), .en(en), .top_left({trees[1394], lumberyards[1394]}), .top({trees[1395], lumberyards[1395]}), .top_right({trees[1396], lumberyards[1396]}), .left({trees[1444], lumberyards[1444]}), .right({trees[1446], lumberyards[1446]}), .bottom_left({trees[1494], lumberyards[1494]}), .bottom({trees[1495], lumberyards[1495]}), .bottom_right({trees[1496], lumberyards[1496]}), .init(2'b00), .state({trees[1445], lumberyards[1445]}));
acre acre_28_46 (.clk(clk), .en(en), .top_left({trees[1395], lumberyards[1395]}), .top({trees[1396], lumberyards[1396]}), .top_right({trees[1397], lumberyards[1397]}), .left({trees[1445], lumberyards[1445]}), .right({trees[1447], lumberyards[1447]}), .bottom_left({trees[1495], lumberyards[1495]}), .bottom({trees[1496], lumberyards[1496]}), .bottom_right({trees[1497], lumberyards[1497]}), .init(2'b10), .state({trees[1446], lumberyards[1446]}));
acre acre_28_47 (.clk(clk), .en(en), .top_left({trees[1396], lumberyards[1396]}), .top({trees[1397], lumberyards[1397]}), .top_right({trees[1398], lumberyards[1398]}), .left({trees[1446], lumberyards[1446]}), .right({trees[1448], lumberyards[1448]}), .bottom_left({trees[1496], lumberyards[1496]}), .bottom({trees[1497], lumberyards[1497]}), .bottom_right({trees[1498], lumberyards[1498]}), .init(2'b00), .state({trees[1447], lumberyards[1447]}));
acre acre_28_48 (.clk(clk), .en(en), .top_left({trees[1397], lumberyards[1397]}), .top({trees[1398], lumberyards[1398]}), .top_right({trees[1399], lumberyards[1399]}), .left({trees[1447], lumberyards[1447]}), .right({trees[1449], lumberyards[1449]}), .bottom_left({trees[1497], lumberyards[1497]}), .bottom({trees[1498], lumberyards[1498]}), .bottom_right({trees[1499], lumberyards[1499]}), .init(2'b00), .state({trees[1448], lumberyards[1448]}));
acre acre_28_49 (.clk(clk), .en(en), .top_left({trees[1398], lumberyards[1398]}), .top({trees[1399], lumberyards[1399]}), .top_right(2'b0), .left({trees[1448], lumberyards[1448]}), .right(2'b0), .bottom_left({trees[1498], lumberyards[1498]}), .bottom({trees[1499], lumberyards[1499]}), .bottom_right(2'b0), .init(2'b00), .state({trees[1449], lumberyards[1449]}));
acre acre_29_0 (.clk(clk), .en(en), .top_left(2'b0), .top({trees[1400], lumberyards[1400]}), .top_right({trees[1401], lumberyards[1401]}), .left(2'b0), .right({trees[1451], lumberyards[1451]}), .bottom_left(2'b0), .bottom({trees[1500], lumberyards[1500]}), .bottom_right({trees[1501], lumberyards[1501]}), .init(2'b00), .state({trees[1450], lumberyards[1450]}));
acre acre_29_1 (.clk(clk), .en(en), .top_left({trees[1400], lumberyards[1400]}), .top({trees[1401], lumberyards[1401]}), .top_right({trees[1402], lumberyards[1402]}), .left({trees[1450], lumberyards[1450]}), .right({trees[1452], lumberyards[1452]}), .bottom_left({trees[1500], lumberyards[1500]}), .bottom({trees[1501], lumberyards[1501]}), .bottom_right({trees[1502], lumberyards[1502]}), .init(2'b10), .state({trees[1451], lumberyards[1451]}));
acre acre_29_2 (.clk(clk), .en(en), .top_left({trees[1401], lumberyards[1401]}), .top({trees[1402], lumberyards[1402]}), .top_right({trees[1403], lumberyards[1403]}), .left({trees[1451], lumberyards[1451]}), .right({trees[1453], lumberyards[1453]}), .bottom_left({trees[1501], lumberyards[1501]}), .bottom({trees[1502], lumberyards[1502]}), .bottom_right({trees[1503], lumberyards[1503]}), .init(2'b10), .state({trees[1452], lumberyards[1452]}));
acre acre_29_3 (.clk(clk), .en(en), .top_left({trees[1402], lumberyards[1402]}), .top({trees[1403], lumberyards[1403]}), .top_right({trees[1404], lumberyards[1404]}), .left({trees[1452], lumberyards[1452]}), .right({trees[1454], lumberyards[1454]}), .bottom_left({trees[1502], lumberyards[1502]}), .bottom({trees[1503], lumberyards[1503]}), .bottom_right({trees[1504], lumberyards[1504]}), .init(2'b00), .state({trees[1453], lumberyards[1453]}));
acre acre_29_4 (.clk(clk), .en(en), .top_left({trees[1403], lumberyards[1403]}), .top({trees[1404], lumberyards[1404]}), .top_right({trees[1405], lumberyards[1405]}), .left({trees[1453], lumberyards[1453]}), .right({trees[1455], lumberyards[1455]}), .bottom_left({trees[1503], lumberyards[1503]}), .bottom({trees[1504], lumberyards[1504]}), .bottom_right({trees[1505], lumberyards[1505]}), .init(2'b00), .state({trees[1454], lumberyards[1454]}));
acre acre_29_5 (.clk(clk), .en(en), .top_left({trees[1404], lumberyards[1404]}), .top({trees[1405], lumberyards[1405]}), .top_right({trees[1406], lumberyards[1406]}), .left({trees[1454], lumberyards[1454]}), .right({trees[1456], lumberyards[1456]}), .bottom_left({trees[1504], lumberyards[1504]}), .bottom({trees[1505], lumberyards[1505]}), .bottom_right({trees[1506], lumberyards[1506]}), .init(2'b00), .state({trees[1455], lumberyards[1455]}));
acre acre_29_6 (.clk(clk), .en(en), .top_left({trees[1405], lumberyards[1405]}), .top({trees[1406], lumberyards[1406]}), .top_right({trees[1407], lumberyards[1407]}), .left({trees[1455], lumberyards[1455]}), .right({trees[1457], lumberyards[1457]}), .bottom_left({trees[1505], lumberyards[1505]}), .bottom({trees[1506], lumberyards[1506]}), .bottom_right({trees[1507], lumberyards[1507]}), .init(2'b00), .state({trees[1456], lumberyards[1456]}));
acre acre_29_7 (.clk(clk), .en(en), .top_left({trees[1406], lumberyards[1406]}), .top({trees[1407], lumberyards[1407]}), .top_right({trees[1408], lumberyards[1408]}), .left({trees[1456], lumberyards[1456]}), .right({trees[1458], lumberyards[1458]}), .bottom_left({trees[1506], lumberyards[1506]}), .bottom({trees[1507], lumberyards[1507]}), .bottom_right({trees[1508], lumberyards[1508]}), .init(2'b01), .state({trees[1457], lumberyards[1457]}));
acre acre_29_8 (.clk(clk), .en(en), .top_left({trees[1407], lumberyards[1407]}), .top({trees[1408], lumberyards[1408]}), .top_right({trees[1409], lumberyards[1409]}), .left({trees[1457], lumberyards[1457]}), .right({trees[1459], lumberyards[1459]}), .bottom_left({trees[1507], lumberyards[1507]}), .bottom({trees[1508], lumberyards[1508]}), .bottom_right({trees[1509], lumberyards[1509]}), .init(2'b00), .state({trees[1458], lumberyards[1458]}));
acre acre_29_9 (.clk(clk), .en(en), .top_left({trees[1408], lumberyards[1408]}), .top({trees[1409], lumberyards[1409]}), .top_right({trees[1410], lumberyards[1410]}), .left({trees[1458], lumberyards[1458]}), .right({trees[1460], lumberyards[1460]}), .bottom_left({trees[1508], lumberyards[1508]}), .bottom({trees[1509], lumberyards[1509]}), .bottom_right({trees[1510], lumberyards[1510]}), .init(2'b00), .state({trees[1459], lumberyards[1459]}));
acre acre_29_10 (.clk(clk), .en(en), .top_left({trees[1409], lumberyards[1409]}), .top({trees[1410], lumberyards[1410]}), .top_right({trees[1411], lumberyards[1411]}), .left({trees[1459], lumberyards[1459]}), .right({trees[1461], lumberyards[1461]}), .bottom_left({trees[1509], lumberyards[1509]}), .bottom({trees[1510], lumberyards[1510]}), .bottom_right({trees[1511], lumberyards[1511]}), .init(2'b10), .state({trees[1460], lumberyards[1460]}));
acre acre_29_11 (.clk(clk), .en(en), .top_left({trees[1410], lumberyards[1410]}), .top({trees[1411], lumberyards[1411]}), .top_right({trees[1412], lumberyards[1412]}), .left({trees[1460], lumberyards[1460]}), .right({trees[1462], lumberyards[1462]}), .bottom_left({trees[1510], lumberyards[1510]}), .bottom({trees[1511], lumberyards[1511]}), .bottom_right({trees[1512], lumberyards[1512]}), .init(2'b10), .state({trees[1461], lumberyards[1461]}));
acre acre_29_12 (.clk(clk), .en(en), .top_left({trees[1411], lumberyards[1411]}), .top({trees[1412], lumberyards[1412]}), .top_right({trees[1413], lumberyards[1413]}), .left({trees[1461], lumberyards[1461]}), .right({trees[1463], lumberyards[1463]}), .bottom_left({trees[1511], lumberyards[1511]}), .bottom({trees[1512], lumberyards[1512]}), .bottom_right({trees[1513], lumberyards[1513]}), .init(2'b10), .state({trees[1462], lumberyards[1462]}));
acre acre_29_13 (.clk(clk), .en(en), .top_left({trees[1412], lumberyards[1412]}), .top({trees[1413], lumberyards[1413]}), .top_right({trees[1414], lumberyards[1414]}), .left({trees[1462], lumberyards[1462]}), .right({trees[1464], lumberyards[1464]}), .bottom_left({trees[1512], lumberyards[1512]}), .bottom({trees[1513], lumberyards[1513]}), .bottom_right({trees[1514], lumberyards[1514]}), .init(2'b00), .state({trees[1463], lumberyards[1463]}));
acre acre_29_14 (.clk(clk), .en(en), .top_left({trees[1413], lumberyards[1413]}), .top({trees[1414], lumberyards[1414]}), .top_right({trees[1415], lumberyards[1415]}), .left({trees[1463], lumberyards[1463]}), .right({trees[1465], lumberyards[1465]}), .bottom_left({trees[1513], lumberyards[1513]}), .bottom({trees[1514], lumberyards[1514]}), .bottom_right({trees[1515], lumberyards[1515]}), .init(2'b10), .state({trees[1464], lumberyards[1464]}));
acre acre_29_15 (.clk(clk), .en(en), .top_left({trees[1414], lumberyards[1414]}), .top({trees[1415], lumberyards[1415]}), .top_right({trees[1416], lumberyards[1416]}), .left({trees[1464], lumberyards[1464]}), .right({trees[1466], lumberyards[1466]}), .bottom_left({trees[1514], lumberyards[1514]}), .bottom({trees[1515], lumberyards[1515]}), .bottom_right({trees[1516], lumberyards[1516]}), .init(2'b01), .state({trees[1465], lumberyards[1465]}));
acre acre_29_16 (.clk(clk), .en(en), .top_left({trees[1415], lumberyards[1415]}), .top({trees[1416], lumberyards[1416]}), .top_right({trees[1417], lumberyards[1417]}), .left({trees[1465], lumberyards[1465]}), .right({trees[1467], lumberyards[1467]}), .bottom_left({trees[1515], lumberyards[1515]}), .bottom({trees[1516], lumberyards[1516]}), .bottom_right({trees[1517], lumberyards[1517]}), .init(2'b00), .state({trees[1466], lumberyards[1466]}));
acre acre_29_17 (.clk(clk), .en(en), .top_left({trees[1416], lumberyards[1416]}), .top({trees[1417], lumberyards[1417]}), .top_right({trees[1418], lumberyards[1418]}), .left({trees[1466], lumberyards[1466]}), .right({trees[1468], lumberyards[1468]}), .bottom_left({trees[1516], lumberyards[1516]}), .bottom({trees[1517], lumberyards[1517]}), .bottom_right({trees[1518], lumberyards[1518]}), .init(2'b00), .state({trees[1467], lumberyards[1467]}));
acre acre_29_18 (.clk(clk), .en(en), .top_left({trees[1417], lumberyards[1417]}), .top({trees[1418], lumberyards[1418]}), .top_right({trees[1419], lumberyards[1419]}), .left({trees[1467], lumberyards[1467]}), .right({trees[1469], lumberyards[1469]}), .bottom_left({trees[1517], lumberyards[1517]}), .bottom({trees[1518], lumberyards[1518]}), .bottom_right({trees[1519], lumberyards[1519]}), .init(2'b01), .state({trees[1468], lumberyards[1468]}));
acre acre_29_19 (.clk(clk), .en(en), .top_left({trees[1418], lumberyards[1418]}), .top({trees[1419], lumberyards[1419]}), .top_right({trees[1420], lumberyards[1420]}), .left({trees[1468], lumberyards[1468]}), .right({trees[1470], lumberyards[1470]}), .bottom_left({trees[1518], lumberyards[1518]}), .bottom({trees[1519], lumberyards[1519]}), .bottom_right({trees[1520], lumberyards[1520]}), .init(2'b00), .state({trees[1469], lumberyards[1469]}));
acre acre_29_20 (.clk(clk), .en(en), .top_left({trees[1419], lumberyards[1419]}), .top({trees[1420], lumberyards[1420]}), .top_right({trees[1421], lumberyards[1421]}), .left({trees[1469], lumberyards[1469]}), .right({trees[1471], lumberyards[1471]}), .bottom_left({trees[1519], lumberyards[1519]}), .bottom({trees[1520], lumberyards[1520]}), .bottom_right({trees[1521], lumberyards[1521]}), .init(2'b00), .state({trees[1470], lumberyards[1470]}));
acre acre_29_21 (.clk(clk), .en(en), .top_left({trees[1420], lumberyards[1420]}), .top({trees[1421], lumberyards[1421]}), .top_right({trees[1422], lumberyards[1422]}), .left({trees[1470], lumberyards[1470]}), .right({trees[1472], lumberyards[1472]}), .bottom_left({trees[1520], lumberyards[1520]}), .bottom({trees[1521], lumberyards[1521]}), .bottom_right({trees[1522], lumberyards[1522]}), .init(2'b00), .state({trees[1471], lumberyards[1471]}));
acre acre_29_22 (.clk(clk), .en(en), .top_left({trees[1421], lumberyards[1421]}), .top({trees[1422], lumberyards[1422]}), .top_right({trees[1423], lumberyards[1423]}), .left({trees[1471], lumberyards[1471]}), .right({trees[1473], lumberyards[1473]}), .bottom_left({trees[1521], lumberyards[1521]}), .bottom({trees[1522], lumberyards[1522]}), .bottom_right({trees[1523], lumberyards[1523]}), .init(2'b00), .state({trees[1472], lumberyards[1472]}));
acre acre_29_23 (.clk(clk), .en(en), .top_left({trees[1422], lumberyards[1422]}), .top({trees[1423], lumberyards[1423]}), .top_right({trees[1424], lumberyards[1424]}), .left({trees[1472], lumberyards[1472]}), .right({trees[1474], lumberyards[1474]}), .bottom_left({trees[1522], lumberyards[1522]}), .bottom({trees[1523], lumberyards[1523]}), .bottom_right({trees[1524], lumberyards[1524]}), .init(2'b00), .state({trees[1473], lumberyards[1473]}));
acre acre_29_24 (.clk(clk), .en(en), .top_left({trees[1423], lumberyards[1423]}), .top({trees[1424], lumberyards[1424]}), .top_right({trees[1425], lumberyards[1425]}), .left({trees[1473], lumberyards[1473]}), .right({trees[1475], lumberyards[1475]}), .bottom_left({trees[1523], lumberyards[1523]}), .bottom({trees[1524], lumberyards[1524]}), .bottom_right({trees[1525], lumberyards[1525]}), .init(2'b00), .state({trees[1474], lumberyards[1474]}));
acre acre_29_25 (.clk(clk), .en(en), .top_left({trees[1424], lumberyards[1424]}), .top({trees[1425], lumberyards[1425]}), .top_right({trees[1426], lumberyards[1426]}), .left({trees[1474], lumberyards[1474]}), .right({trees[1476], lumberyards[1476]}), .bottom_left({trees[1524], lumberyards[1524]}), .bottom({trees[1525], lumberyards[1525]}), .bottom_right({trees[1526], lumberyards[1526]}), .init(2'b10), .state({trees[1475], lumberyards[1475]}));
acre acre_29_26 (.clk(clk), .en(en), .top_left({trees[1425], lumberyards[1425]}), .top({trees[1426], lumberyards[1426]}), .top_right({trees[1427], lumberyards[1427]}), .left({trees[1475], lumberyards[1475]}), .right({trees[1477], lumberyards[1477]}), .bottom_left({trees[1525], lumberyards[1525]}), .bottom({trees[1526], lumberyards[1526]}), .bottom_right({trees[1527], lumberyards[1527]}), .init(2'b10), .state({trees[1476], lumberyards[1476]}));
acre acre_29_27 (.clk(clk), .en(en), .top_left({trees[1426], lumberyards[1426]}), .top({trees[1427], lumberyards[1427]}), .top_right({trees[1428], lumberyards[1428]}), .left({trees[1476], lumberyards[1476]}), .right({trees[1478], lumberyards[1478]}), .bottom_left({trees[1526], lumberyards[1526]}), .bottom({trees[1527], lumberyards[1527]}), .bottom_right({trees[1528], lumberyards[1528]}), .init(2'b10), .state({trees[1477], lumberyards[1477]}));
acre acre_29_28 (.clk(clk), .en(en), .top_left({trees[1427], lumberyards[1427]}), .top({trees[1428], lumberyards[1428]}), .top_right({trees[1429], lumberyards[1429]}), .left({trees[1477], lumberyards[1477]}), .right({trees[1479], lumberyards[1479]}), .bottom_left({trees[1527], lumberyards[1527]}), .bottom({trees[1528], lumberyards[1528]}), .bottom_right({trees[1529], lumberyards[1529]}), .init(2'b00), .state({trees[1478], lumberyards[1478]}));
acre acre_29_29 (.clk(clk), .en(en), .top_left({trees[1428], lumberyards[1428]}), .top({trees[1429], lumberyards[1429]}), .top_right({trees[1430], lumberyards[1430]}), .left({trees[1478], lumberyards[1478]}), .right({trees[1480], lumberyards[1480]}), .bottom_left({trees[1528], lumberyards[1528]}), .bottom({trees[1529], lumberyards[1529]}), .bottom_right({trees[1530], lumberyards[1530]}), .init(2'b00), .state({trees[1479], lumberyards[1479]}));
acre acre_29_30 (.clk(clk), .en(en), .top_left({trees[1429], lumberyards[1429]}), .top({trees[1430], lumberyards[1430]}), .top_right({trees[1431], lumberyards[1431]}), .left({trees[1479], lumberyards[1479]}), .right({trees[1481], lumberyards[1481]}), .bottom_left({trees[1529], lumberyards[1529]}), .bottom({trees[1530], lumberyards[1530]}), .bottom_right({trees[1531], lumberyards[1531]}), .init(2'b00), .state({trees[1480], lumberyards[1480]}));
acre acre_29_31 (.clk(clk), .en(en), .top_left({trees[1430], lumberyards[1430]}), .top({trees[1431], lumberyards[1431]}), .top_right({trees[1432], lumberyards[1432]}), .left({trees[1480], lumberyards[1480]}), .right({trees[1482], lumberyards[1482]}), .bottom_left({trees[1530], lumberyards[1530]}), .bottom({trees[1531], lumberyards[1531]}), .bottom_right({trees[1532], lumberyards[1532]}), .init(2'b00), .state({trees[1481], lumberyards[1481]}));
acre acre_29_32 (.clk(clk), .en(en), .top_left({trees[1431], lumberyards[1431]}), .top({trees[1432], lumberyards[1432]}), .top_right({trees[1433], lumberyards[1433]}), .left({trees[1481], lumberyards[1481]}), .right({trees[1483], lumberyards[1483]}), .bottom_left({trees[1531], lumberyards[1531]}), .bottom({trees[1532], lumberyards[1532]}), .bottom_right({trees[1533], lumberyards[1533]}), .init(2'b10), .state({trees[1482], lumberyards[1482]}));
acre acre_29_33 (.clk(clk), .en(en), .top_left({trees[1432], lumberyards[1432]}), .top({trees[1433], lumberyards[1433]}), .top_right({trees[1434], lumberyards[1434]}), .left({trees[1482], lumberyards[1482]}), .right({trees[1484], lumberyards[1484]}), .bottom_left({trees[1532], lumberyards[1532]}), .bottom({trees[1533], lumberyards[1533]}), .bottom_right({trees[1534], lumberyards[1534]}), .init(2'b00), .state({trees[1483], lumberyards[1483]}));
acre acre_29_34 (.clk(clk), .en(en), .top_left({trees[1433], lumberyards[1433]}), .top({trees[1434], lumberyards[1434]}), .top_right({trees[1435], lumberyards[1435]}), .left({trees[1483], lumberyards[1483]}), .right({trees[1485], lumberyards[1485]}), .bottom_left({trees[1533], lumberyards[1533]}), .bottom({trees[1534], lumberyards[1534]}), .bottom_right({trees[1535], lumberyards[1535]}), .init(2'b00), .state({trees[1484], lumberyards[1484]}));
acre acre_29_35 (.clk(clk), .en(en), .top_left({trees[1434], lumberyards[1434]}), .top({trees[1435], lumberyards[1435]}), .top_right({trees[1436], lumberyards[1436]}), .left({trees[1484], lumberyards[1484]}), .right({trees[1486], lumberyards[1486]}), .bottom_left({trees[1534], lumberyards[1534]}), .bottom({trees[1535], lumberyards[1535]}), .bottom_right({trees[1536], lumberyards[1536]}), .init(2'b00), .state({trees[1485], lumberyards[1485]}));
acre acre_29_36 (.clk(clk), .en(en), .top_left({trees[1435], lumberyards[1435]}), .top({trees[1436], lumberyards[1436]}), .top_right({trees[1437], lumberyards[1437]}), .left({trees[1485], lumberyards[1485]}), .right({trees[1487], lumberyards[1487]}), .bottom_left({trees[1535], lumberyards[1535]}), .bottom({trees[1536], lumberyards[1536]}), .bottom_right({trees[1537], lumberyards[1537]}), .init(2'b01), .state({trees[1486], lumberyards[1486]}));
acre acre_29_37 (.clk(clk), .en(en), .top_left({trees[1436], lumberyards[1436]}), .top({trees[1437], lumberyards[1437]}), .top_right({trees[1438], lumberyards[1438]}), .left({trees[1486], lumberyards[1486]}), .right({trees[1488], lumberyards[1488]}), .bottom_left({trees[1536], lumberyards[1536]}), .bottom({trees[1537], lumberyards[1537]}), .bottom_right({trees[1538], lumberyards[1538]}), .init(2'b00), .state({trees[1487], lumberyards[1487]}));
acre acre_29_38 (.clk(clk), .en(en), .top_left({trees[1437], lumberyards[1437]}), .top({trees[1438], lumberyards[1438]}), .top_right({trees[1439], lumberyards[1439]}), .left({trees[1487], lumberyards[1487]}), .right({trees[1489], lumberyards[1489]}), .bottom_left({trees[1537], lumberyards[1537]}), .bottom({trees[1538], lumberyards[1538]}), .bottom_right({trees[1539], lumberyards[1539]}), .init(2'b00), .state({trees[1488], lumberyards[1488]}));
acre acre_29_39 (.clk(clk), .en(en), .top_left({trees[1438], lumberyards[1438]}), .top({trees[1439], lumberyards[1439]}), .top_right({trees[1440], lumberyards[1440]}), .left({trees[1488], lumberyards[1488]}), .right({trees[1490], lumberyards[1490]}), .bottom_left({trees[1538], lumberyards[1538]}), .bottom({trees[1539], lumberyards[1539]}), .bottom_right({trees[1540], lumberyards[1540]}), .init(2'b01), .state({trees[1489], lumberyards[1489]}));
acre acre_29_40 (.clk(clk), .en(en), .top_left({trees[1439], lumberyards[1439]}), .top({trees[1440], lumberyards[1440]}), .top_right({trees[1441], lumberyards[1441]}), .left({trees[1489], lumberyards[1489]}), .right({trees[1491], lumberyards[1491]}), .bottom_left({trees[1539], lumberyards[1539]}), .bottom({trees[1540], lumberyards[1540]}), .bottom_right({trees[1541], lumberyards[1541]}), .init(2'b00), .state({trees[1490], lumberyards[1490]}));
acre acre_29_41 (.clk(clk), .en(en), .top_left({trees[1440], lumberyards[1440]}), .top({trees[1441], lumberyards[1441]}), .top_right({trees[1442], lumberyards[1442]}), .left({trees[1490], lumberyards[1490]}), .right({trees[1492], lumberyards[1492]}), .bottom_left({trees[1540], lumberyards[1540]}), .bottom({trees[1541], lumberyards[1541]}), .bottom_right({trees[1542], lumberyards[1542]}), .init(2'b10), .state({trees[1491], lumberyards[1491]}));
acre acre_29_42 (.clk(clk), .en(en), .top_left({trees[1441], lumberyards[1441]}), .top({trees[1442], lumberyards[1442]}), .top_right({trees[1443], lumberyards[1443]}), .left({trees[1491], lumberyards[1491]}), .right({trees[1493], lumberyards[1493]}), .bottom_left({trees[1541], lumberyards[1541]}), .bottom({trees[1542], lumberyards[1542]}), .bottom_right({trees[1543], lumberyards[1543]}), .init(2'b10), .state({trees[1492], lumberyards[1492]}));
acre acre_29_43 (.clk(clk), .en(en), .top_left({trees[1442], lumberyards[1442]}), .top({trees[1443], lumberyards[1443]}), .top_right({trees[1444], lumberyards[1444]}), .left({trees[1492], lumberyards[1492]}), .right({trees[1494], lumberyards[1494]}), .bottom_left({trees[1542], lumberyards[1542]}), .bottom({trees[1543], lumberyards[1543]}), .bottom_right({trees[1544], lumberyards[1544]}), .init(2'b00), .state({trees[1493], lumberyards[1493]}));
acre acre_29_44 (.clk(clk), .en(en), .top_left({trees[1443], lumberyards[1443]}), .top({trees[1444], lumberyards[1444]}), .top_right({trees[1445], lumberyards[1445]}), .left({trees[1493], lumberyards[1493]}), .right({trees[1495], lumberyards[1495]}), .bottom_left({trees[1543], lumberyards[1543]}), .bottom({trees[1544], lumberyards[1544]}), .bottom_right({trees[1545], lumberyards[1545]}), .init(2'b00), .state({trees[1494], lumberyards[1494]}));
acre acre_29_45 (.clk(clk), .en(en), .top_left({trees[1444], lumberyards[1444]}), .top({trees[1445], lumberyards[1445]}), .top_right({trees[1446], lumberyards[1446]}), .left({trees[1494], lumberyards[1494]}), .right({trees[1496], lumberyards[1496]}), .bottom_left({trees[1544], lumberyards[1544]}), .bottom({trees[1545], lumberyards[1545]}), .bottom_right({trees[1546], lumberyards[1546]}), .init(2'b10), .state({trees[1495], lumberyards[1495]}));
acre acre_29_46 (.clk(clk), .en(en), .top_left({trees[1445], lumberyards[1445]}), .top({trees[1446], lumberyards[1446]}), .top_right({trees[1447], lumberyards[1447]}), .left({trees[1495], lumberyards[1495]}), .right({trees[1497], lumberyards[1497]}), .bottom_left({trees[1545], lumberyards[1545]}), .bottom({trees[1546], lumberyards[1546]}), .bottom_right({trees[1547], lumberyards[1547]}), .init(2'b00), .state({trees[1496], lumberyards[1496]}));
acre acre_29_47 (.clk(clk), .en(en), .top_left({trees[1446], lumberyards[1446]}), .top({trees[1447], lumberyards[1447]}), .top_right({trees[1448], lumberyards[1448]}), .left({trees[1496], lumberyards[1496]}), .right({trees[1498], lumberyards[1498]}), .bottom_left({trees[1546], lumberyards[1546]}), .bottom({trees[1547], lumberyards[1547]}), .bottom_right({trees[1548], lumberyards[1548]}), .init(2'b00), .state({trees[1497], lumberyards[1497]}));
acre acre_29_48 (.clk(clk), .en(en), .top_left({trees[1447], lumberyards[1447]}), .top({trees[1448], lumberyards[1448]}), .top_right({trees[1449], lumberyards[1449]}), .left({trees[1497], lumberyards[1497]}), .right({trees[1499], lumberyards[1499]}), .bottom_left({trees[1547], lumberyards[1547]}), .bottom({trees[1548], lumberyards[1548]}), .bottom_right({trees[1549], lumberyards[1549]}), .init(2'b00), .state({trees[1498], lumberyards[1498]}));
acre acre_29_49 (.clk(clk), .en(en), .top_left({trees[1448], lumberyards[1448]}), .top({trees[1449], lumberyards[1449]}), .top_right(2'b0), .left({trees[1498], lumberyards[1498]}), .right(2'b0), .bottom_left({trees[1548], lumberyards[1548]}), .bottom({trees[1549], lumberyards[1549]}), .bottom_right(2'b0), .init(2'b00), .state({trees[1499], lumberyards[1499]}));
acre acre_30_0 (.clk(clk), .en(en), .top_left(2'b0), .top({trees[1450], lumberyards[1450]}), .top_right({trees[1451], lumberyards[1451]}), .left(2'b0), .right({trees[1501], lumberyards[1501]}), .bottom_left(2'b0), .bottom({trees[1550], lumberyards[1550]}), .bottom_right({trees[1551], lumberyards[1551]}), .init(2'b01), .state({trees[1500], lumberyards[1500]}));
acre acre_30_1 (.clk(clk), .en(en), .top_left({trees[1450], lumberyards[1450]}), .top({trees[1451], lumberyards[1451]}), .top_right({trees[1452], lumberyards[1452]}), .left({trees[1500], lumberyards[1500]}), .right({trees[1502], lumberyards[1502]}), .bottom_left({trees[1550], lumberyards[1550]}), .bottom({trees[1551], lumberyards[1551]}), .bottom_right({trees[1552], lumberyards[1552]}), .init(2'b00), .state({trees[1501], lumberyards[1501]}));
acre acre_30_2 (.clk(clk), .en(en), .top_left({trees[1451], lumberyards[1451]}), .top({trees[1452], lumberyards[1452]}), .top_right({trees[1453], lumberyards[1453]}), .left({trees[1501], lumberyards[1501]}), .right({trees[1503], lumberyards[1503]}), .bottom_left({trees[1551], lumberyards[1551]}), .bottom({trees[1552], lumberyards[1552]}), .bottom_right({trees[1553], lumberyards[1553]}), .init(2'b10), .state({trees[1502], lumberyards[1502]}));
acre acre_30_3 (.clk(clk), .en(en), .top_left({trees[1452], lumberyards[1452]}), .top({trees[1453], lumberyards[1453]}), .top_right({trees[1454], lumberyards[1454]}), .left({trees[1502], lumberyards[1502]}), .right({trees[1504], lumberyards[1504]}), .bottom_left({trees[1552], lumberyards[1552]}), .bottom({trees[1553], lumberyards[1553]}), .bottom_right({trees[1554], lumberyards[1554]}), .init(2'b10), .state({trees[1503], lumberyards[1503]}));
acre acre_30_4 (.clk(clk), .en(en), .top_left({trees[1453], lumberyards[1453]}), .top({trees[1454], lumberyards[1454]}), .top_right({trees[1455], lumberyards[1455]}), .left({trees[1503], lumberyards[1503]}), .right({trees[1505], lumberyards[1505]}), .bottom_left({trees[1553], lumberyards[1553]}), .bottom({trees[1554], lumberyards[1554]}), .bottom_right({trees[1555], lumberyards[1555]}), .init(2'b00), .state({trees[1504], lumberyards[1504]}));
acre acre_30_5 (.clk(clk), .en(en), .top_left({trees[1454], lumberyards[1454]}), .top({trees[1455], lumberyards[1455]}), .top_right({trees[1456], lumberyards[1456]}), .left({trees[1504], lumberyards[1504]}), .right({trees[1506], lumberyards[1506]}), .bottom_left({trees[1554], lumberyards[1554]}), .bottom({trees[1555], lumberyards[1555]}), .bottom_right({trees[1556], lumberyards[1556]}), .init(2'b10), .state({trees[1505], lumberyards[1505]}));
acre acre_30_6 (.clk(clk), .en(en), .top_left({trees[1455], lumberyards[1455]}), .top({trees[1456], lumberyards[1456]}), .top_right({trees[1457], lumberyards[1457]}), .left({trees[1505], lumberyards[1505]}), .right({trees[1507], lumberyards[1507]}), .bottom_left({trees[1555], lumberyards[1555]}), .bottom({trees[1556], lumberyards[1556]}), .bottom_right({trees[1557], lumberyards[1557]}), .init(2'b00), .state({trees[1506], lumberyards[1506]}));
acre acre_30_7 (.clk(clk), .en(en), .top_left({trees[1456], lumberyards[1456]}), .top({trees[1457], lumberyards[1457]}), .top_right({trees[1458], lumberyards[1458]}), .left({trees[1506], lumberyards[1506]}), .right({trees[1508], lumberyards[1508]}), .bottom_left({trees[1556], lumberyards[1556]}), .bottom({trees[1557], lumberyards[1557]}), .bottom_right({trees[1558], lumberyards[1558]}), .init(2'b00), .state({trees[1507], lumberyards[1507]}));
acre acre_30_8 (.clk(clk), .en(en), .top_left({trees[1457], lumberyards[1457]}), .top({trees[1458], lumberyards[1458]}), .top_right({trees[1459], lumberyards[1459]}), .left({trees[1507], lumberyards[1507]}), .right({trees[1509], lumberyards[1509]}), .bottom_left({trees[1557], lumberyards[1557]}), .bottom({trees[1558], lumberyards[1558]}), .bottom_right({trees[1559], lumberyards[1559]}), .init(2'b00), .state({trees[1508], lumberyards[1508]}));
acre acre_30_9 (.clk(clk), .en(en), .top_left({trees[1458], lumberyards[1458]}), .top({trees[1459], lumberyards[1459]}), .top_right({trees[1460], lumberyards[1460]}), .left({trees[1508], lumberyards[1508]}), .right({trees[1510], lumberyards[1510]}), .bottom_left({trees[1558], lumberyards[1558]}), .bottom({trees[1559], lumberyards[1559]}), .bottom_right({trees[1560], lumberyards[1560]}), .init(2'b00), .state({trees[1509], lumberyards[1509]}));
acre acre_30_10 (.clk(clk), .en(en), .top_left({trees[1459], lumberyards[1459]}), .top({trees[1460], lumberyards[1460]}), .top_right({trees[1461], lumberyards[1461]}), .left({trees[1509], lumberyards[1509]}), .right({trees[1511], lumberyards[1511]}), .bottom_left({trees[1559], lumberyards[1559]}), .bottom({trees[1560], lumberyards[1560]}), .bottom_right({trees[1561], lumberyards[1561]}), .init(2'b10), .state({trees[1510], lumberyards[1510]}));
acre acre_30_11 (.clk(clk), .en(en), .top_left({trees[1460], lumberyards[1460]}), .top({trees[1461], lumberyards[1461]}), .top_right({trees[1462], lumberyards[1462]}), .left({trees[1510], lumberyards[1510]}), .right({trees[1512], lumberyards[1512]}), .bottom_left({trees[1560], lumberyards[1560]}), .bottom({trees[1561], lumberyards[1561]}), .bottom_right({trees[1562], lumberyards[1562]}), .init(2'b00), .state({trees[1511], lumberyards[1511]}));
acre acre_30_12 (.clk(clk), .en(en), .top_left({trees[1461], lumberyards[1461]}), .top({trees[1462], lumberyards[1462]}), .top_right({trees[1463], lumberyards[1463]}), .left({trees[1511], lumberyards[1511]}), .right({trees[1513], lumberyards[1513]}), .bottom_left({trees[1561], lumberyards[1561]}), .bottom({trees[1562], lumberyards[1562]}), .bottom_right({trees[1563], lumberyards[1563]}), .init(2'b00), .state({trees[1512], lumberyards[1512]}));
acre acre_30_13 (.clk(clk), .en(en), .top_left({trees[1462], lumberyards[1462]}), .top({trees[1463], lumberyards[1463]}), .top_right({trees[1464], lumberyards[1464]}), .left({trees[1512], lumberyards[1512]}), .right({trees[1514], lumberyards[1514]}), .bottom_left({trees[1562], lumberyards[1562]}), .bottom({trees[1563], lumberyards[1563]}), .bottom_right({trees[1564], lumberyards[1564]}), .init(2'b00), .state({trees[1513], lumberyards[1513]}));
acre acre_30_14 (.clk(clk), .en(en), .top_left({trees[1463], lumberyards[1463]}), .top({trees[1464], lumberyards[1464]}), .top_right({trees[1465], lumberyards[1465]}), .left({trees[1513], lumberyards[1513]}), .right({trees[1515], lumberyards[1515]}), .bottom_left({trees[1563], lumberyards[1563]}), .bottom({trees[1564], lumberyards[1564]}), .bottom_right({trees[1565], lumberyards[1565]}), .init(2'b00), .state({trees[1514], lumberyards[1514]}));
acre acre_30_15 (.clk(clk), .en(en), .top_left({trees[1464], lumberyards[1464]}), .top({trees[1465], lumberyards[1465]}), .top_right({trees[1466], lumberyards[1466]}), .left({trees[1514], lumberyards[1514]}), .right({trees[1516], lumberyards[1516]}), .bottom_left({trees[1564], lumberyards[1564]}), .bottom({trees[1565], lumberyards[1565]}), .bottom_right({trees[1566], lumberyards[1566]}), .init(2'b00), .state({trees[1515], lumberyards[1515]}));
acre acre_30_16 (.clk(clk), .en(en), .top_left({trees[1465], lumberyards[1465]}), .top({trees[1466], lumberyards[1466]}), .top_right({trees[1467], lumberyards[1467]}), .left({trees[1515], lumberyards[1515]}), .right({trees[1517], lumberyards[1517]}), .bottom_left({trees[1565], lumberyards[1565]}), .bottom({trees[1566], lumberyards[1566]}), .bottom_right({trees[1567], lumberyards[1567]}), .init(2'b00), .state({trees[1516], lumberyards[1516]}));
acre acre_30_17 (.clk(clk), .en(en), .top_left({trees[1466], lumberyards[1466]}), .top({trees[1467], lumberyards[1467]}), .top_right({trees[1468], lumberyards[1468]}), .left({trees[1516], lumberyards[1516]}), .right({trees[1518], lumberyards[1518]}), .bottom_left({trees[1566], lumberyards[1566]}), .bottom({trees[1567], lumberyards[1567]}), .bottom_right({trees[1568], lumberyards[1568]}), .init(2'b00), .state({trees[1517], lumberyards[1517]}));
acre acre_30_18 (.clk(clk), .en(en), .top_left({trees[1467], lumberyards[1467]}), .top({trees[1468], lumberyards[1468]}), .top_right({trees[1469], lumberyards[1469]}), .left({trees[1517], lumberyards[1517]}), .right({trees[1519], lumberyards[1519]}), .bottom_left({trees[1567], lumberyards[1567]}), .bottom({trees[1568], lumberyards[1568]}), .bottom_right({trees[1569], lumberyards[1569]}), .init(2'b00), .state({trees[1518], lumberyards[1518]}));
acre acre_30_19 (.clk(clk), .en(en), .top_left({trees[1468], lumberyards[1468]}), .top({trees[1469], lumberyards[1469]}), .top_right({trees[1470], lumberyards[1470]}), .left({trees[1518], lumberyards[1518]}), .right({trees[1520], lumberyards[1520]}), .bottom_left({trees[1568], lumberyards[1568]}), .bottom({trees[1569], lumberyards[1569]}), .bottom_right({trees[1570], lumberyards[1570]}), .init(2'b00), .state({trees[1519], lumberyards[1519]}));
acre acre_30_20 (.clk(clk), .en(en), .top_left({trees[1469], lumberyards[1469]}), .top({trees[1470], lumberyards[1470]}), .top_right({trees[1471], lumberyards[1471]}), .left({trees[1519], lumberyards[1519]}), .right({trees[1521], lumberyards[1521]}), .bottom_left({trees[1569], lumberyards[1569]}), .bottom({trees[1570], lumberyards[1570]}), .bottom_right({trees[1571], lumberyards[1571]}), .init(2'b00), .state({trees[1520], lumberyards[1520]}));
acre acre_30_21 (.clk(clk), .en(en), .top_left({trees[1470], lumberyards[1470]}), .top({trees[1471], lumberyards[1471]}), .top_right({trees[1472], lumberyards[1472]}), .left({trees[1520], lumberyards[1520]}), .right({trees[1522], lumberyards[1522]}), .bottom_left({trees[1570], lumberyards[1570]}), .bottom({trees[1571], lumberyards[1571]}), .bottom_right({trees[1572], lumberyards[1572]}), .init(2'b10), .state({trees[1521], lumberyards[1521]}));
acre acre_30_22 (.clk(clk), .en(en), .top_left({trees[1471], lumberyards[1471]}), .top({trees[1472], lumberyards[1472]}), .top_right({trees[1473], lumberyards[1473]}), .left({trees[1521], lumberyards[1521]}), .right({trees[1523], lumberyards[1523]}), .bottom_left({trees[1571], lumberyards[1571]}), .bottom({trees[1572], lumberyards[1572]}), .bottom_right({trees[1573], lumberyards[1573]}), .init(2'b00), .state({trees[1522], lumberyards[1522]}));
acre acre_30_23 (.clk(clk), .en(en), .top_left({trees[1472], lumberyards[1472]}), .top({trees[1473], lumberyards[1473]}), .top_right({trees[1474], lumberyards[1474]}), .left({trees[1522], lumberyards[1522]}), .right({trees[1524], lumberyards[1524]}), .bottom_left({trees[1572], lumberyards[1572]}), .bottom({trees[1573], lumberyards[1573]}), .bottom_right({trees[1574], lumberyards[1574]}), .init(2'b10), .state({trees[1523], lumberyards[1523]}));
acre acre_30_24 (.clk(clk), .en(en), .top_left({trees[1473], lumberyards[1473]}), .top({trees[1474], lumberyards[1474]}), .top_right({trees[1475], lumberyards[1475]}), .left({trees[1523], lumberyards[1523]}), .right({trees[1525], lumberyards[1525]}), .bottom_left({trees[1573], lumberyards[1573]}), .bottom({trees[1574], lumberyards[1574]}), .bottom_right({trees[1575], lumberyards[1575]}), .init(2'b00), .state({trees[1524], lumberyards[1524]}));
acre acre_30_25 (.clk(clk), .en(en), .top_left({trees[1474], lumberyards[1474]}), .top({trees[1475], lumberyards[1475]}), .top_right({trees[1476], lumberyards[1476]}), .left({trees[1524], lumberyards[1524]}), .right({trees[1526], lumberyards[1526]}), .bottom_left({trees[1574], lumberyards[1574]}), .bottom({trees[1575], lumberyards[1575]}), .bottom_right({trees[1576], lumberyards[1576]}), .init(2'b00), .state({trees[1525], lumberyards[1525]}));
acre acre_30_26 (.clk(clk), .en(en), .top_left({trees[1475], lumberyards[1475]}), .top({trees[1476], lumberyards[1476]}), .top_right({trees[1477], lumberyards[1477]}), .left({trees[1525], lumberyards[1525]}), .right({trees[1527], lumberyards[1527]}), .bottom_left({trees[1575], lumberyards[1575]}), .bottom({trees[1576], lumberyards[1576]}), .bottom_right({trees[1577], lumberyards[1577]}), .init(2'b00), .state({trees[1526], lumberyards[1526]}));
acre acre_30_27 (.clk(clk), .en(en), .top_left({trees[1476], lumberyards[1476]}), .top({trees[1477], lumberyards[1477]}), .top_right({trees[1478], lumberyards[1478]}), .left({trees[1526], lumberyards[1526]}), .right({trees[1528], lumberyards[1528]}), .bottom_left({trees[1576], lumberyards[1576]}), .bottom({trees[1577], lumberyards[1577]}), .bottom_right({trees[1578], lumberyards[1578]}), .init(2'b01), .state({trees[1527], lumberyards[1527]}));
acre acre_30_28 (.clk(clk), .en(en), .top_left({trees[1477], lumberyards[1477]}), .top({trees[1478], lumberyards[1478]}), .top_right({trees[1479], lumberyards[1479]}), .left({trees[1527], lumberyards[1527]}), .right({trees[1529], lumberyards[1529]}), .bottom_left({trees[1577], lumberyards[1577]}), .bottom({trees[1578], lumberyards[1578]}), .bottom_right({trees[1579], lumberyards[1579]}), .init(2'b01), .state({trees[1528], lumberyards[1528]}));
acre acre_30_29 (.clk(clk), .en(en), .top_left({trees[1478], lumberyards[1478]}), .top({trees[1479], lumberyards[1479]}), .top_right({trees[1480], lumberyards[1480]}), .left({trees[1528], lumberyards[1528]}), .right({trees[1530], lumberyards[1530]}), .bottom_left({trees[1578], lumberyards[1578]}), .bottom({trees[1579], lumberyards[1579]}), .bottom_right({trees[1580], lumberyards[1580]}), .init(2'b10), .state({trees[1529], lumberyards[1529]}));
acre acre_30_30 (.clk(clk), .en(en), .top_left({trees[1479], lumberyards[1479]}), .top({trees[1480], lumberyards[1480]}), .top_right({trees[1481], lumberyards[1481]}), .left({trees[1529], lumberyards[1529]}), .right({trees[1531], lumberyards[1531]}), .bottom_left({trees[1579], lumberyards[1579]}), .bottom({trees[1580], lumberyards[1580]}), .bottom_right({trees[1581], lumberyards[1581]}), .init(2'b01), .state({trees[1530], lumberyards[1530]}));
acre acre_30_31 (.clk(clk), .en(en), .top_left({trees[1480], lumberyards[1480]}), .top({trees[1481], lumberyards[1481]}), .top_right({trees[1482], lumberyards[1482]}), .left({trees[1530], lumberyards[1530]}), .right({trees[1532], lumberyards[1532]}), .bottom_left({trees[1580], lumberyards[1580]}), .bottom({trees[1581], lumberyards[1581]}), .bottom_right({trees[1582], lumberyards[1582]}), .init(2'b10), .state({trees[1531], lumberyards[1531]}));
acre acre_30_32 (.clk(clk), .en(en), .top_left({trees[1481], lumberyards[1481]}), .top({trees[1482], lumberyards[1482]}), .top_right({trees[1483], lumberyards[1483]}), .left({trees[1531], lumberyards[1531]}), .right({trees[1533], lumberyards[1533]}), .bottom_left({trees[1581], lumberyards[1581]}), .bottom({trees[1582], lumberyards[1582]}), .bottom_right({trees[1583], lumberyards[1583]}), .init(2'b00), .state({trees[1532], lumberyards[1532]}));
acre acre_30_33 (.clk(clk), .en(en), .top_left({trees[1482], lumberyards[1482]}), .top({trees[1483], lumberyards[1483]}), .top_right({trees[1484], lumberyards[1484]}), .left({trees[1532], lumberyards[1532]}), .right({trees[1534], lumberyards[1534]}), .bottom_left({trees[1582], lumberyards[1582]}), .bottom({trees[1583], lumberyards[1583]}), .bottom_right({trees[1584], lumberyards[1584]}), .init(2'b00), .state({trees[1533], lumberyards[1533]}));
acre acre_30_34 (.clk(clk), .en(en), .top_left({trees[1483], lumberyards[1483]}), .top({trees[1484], lumberyards[1484]}), .top_right({trees[1485], lumberyards[1485]}), .left({trees[1533], lumberyards[1533]}), .right({trees[1535], lumberyards[1535]}), .bottom_left({trees[1583], lumberyards[1583]}), .bottom({trees[1584], lumberyards[1584]}), .bottom_right({trees[1585], lumberyards[1585]}), .init(2'b10), .state({trees[1534], lumberyards[1534]}));
acre acre_30_35 (.clk(clk), .en(en), .top_left({trees[1484], lumberyards[1484]}), .top({trees[1485], lumberyards[1485]}), .top_right({trees[1486], lumberyards[1486]}), .left({trees[1534], lumberyards[1534]}), .right({trees[1536], lumberyards[1536]}), .bottom_left({trees[1584], lumberyards[1584]}), .bottom({trees[1585], lumberyards[1585]}), .bottom_right({trees[1586], lumberyards[1586]}), .init(2'b01), .state({trees[1535], lumberyards[1535]}));
acre acre_30_36 (.clk(clk), .en(en), .top_left({trees[1485], lumberyards[1485]}), .top({trees[1486], lumberyards[1486]}), .top_right({trees[1487], lumberyards[1487]}), .left({trees[1535], lumberyards[1535]}), .right({trees[1537], lumberyards[1537]}), .bottom_left({trees[1585], lumberyards[1585]}), .bottom({trees[1586], lumberyards[1586]}), .bottom_right({trees[1587], lumberyards[1587]}), .init(2'b00), .state({trees[1536], lumberyards[1536]}));
acre acre_30_37 (.clk(clk), .en(en), .top_left({trees[1486], lumberyards[1486]}), .top({trees[1487], lumberyards[1487]}), .top_right({trees[1488], lumberyards[1488]}), .left({trees[1536], lumberyards[1536]}), .right({trees[1538], lumberyards[1538]}), .bottom_left({trees[1586], lumberyards[1586]}), .bottom({trees[1587], lumberyards[1587]}), .bottom_right({trees[1588], lumberyards[1588]}), .init(2'b00), .state({trees[1537], lumberyards[1537]}));
acre acre_30_38 (.clk(clk), .en(en), .top_left({trees[1487], lumberyards[1487]}), .top({trees[1488], lumberyards[1488]}), .top_right({trees[1489], lumberyards[1489]}), .left({trees[1537], lumberyards[1537]}), .right({trees[1539], lumberyards[1539]}), .bottom_left({trees[1587], lumberyards[1587]}), .bottom({trees[1588], lumberyards[1588]}), .bottom_right({trees[1589], lumberyards[1589]}), .init(2'b00), .state({trees[1538], lumberyards[1538]}));
acre acre_30_39 (.clk(clk), .en(en), .top_left({trees[1488], lumberyards[1488]}), .top({trees[1489], lumberyards[1489]}), .top_right({trees[1490], lumberyards[1490]}), .left({trees[1538], lumberyards[1538]}), .right({trees[1540], lumberyards[1540]}), .bottom_left({trees[1588], lumberyards[1588]}), .bottom({trees[1589], lumberyards[1589]}), .bottom_right({trees[1590], lumberyards[1590]}), .init(2'b00), .state({trees[1539], lumberyards[1539]}));
acre acre_30_40 (.clk(clk), .en(en), .top_left({trees[1489], lumberyards[1489]}), .top({trees[1490], lumberyards[1490]}), .top_right({trees[1491], lumberyards[1491]}), .left({trees[1539], lumberyards[1539]}), .right({trees[1541], lumberyards[1541]}), .bottom_left({trees[1589], lumberyards[1589]}), .bottom({trees[1590], lumberyards[1590]}), .bottom_right({trees[1591], lumberyards[1591]}), .init(2'b10), .state({trees[1540], lumberyards[1540]}));
acre acre_30_41 (.clk(clk), .en(en), .top_left({trees[1490], lumberyards[1490]}), .top({trees[1491], lumberyards[1491]}), .top_right({trees[1492], lumberyards[1492]}), .left({trees[1540], lumberyards[1540]}), .right({trees[1542], lumberyards[1542]}), .bottom_left({trees[1590], lumberyards[1590]}), .bottom({trees[1591], lumberyards[1591]}), .bottom_right({trees[1592], lumberyards[1592]}), .init(2'b00), .state({trees[1541], lumberyards[1541]}));
acre acre_30_42 (.clk(clk), .en(en), .top_left({trees[1491], lumberyards[1491]}), .top({trees[1492], lumberyards[1492]}), .top_right({trees[1493], lumberyards[1493]}), .left({trees[1541], lumberyards[1541]}), .right({trees[1543], lumberyards[1543]}), .bottom_left({trees[1591], lumberyards[1591]}), .bottom({trees[1592], lumberyards[1592]}), .bottom_right({trees[1593], lumberyards[1593]}), .init(2'b01), .state({trees[1542], lumberyards[1542]}));
acre acre_30_43 (.clk(clk), .en(en), .top_left({trees[1492], lumberyards[1492]}), .top({trees[1493], lumberyards[1493]}), .top_right({trees[1494], lumberyards[1494]}), .left({trees[1542], lumberyards[1542]}), .right({trees[1544], lumberyards[1544]}), .bottom_left({trees[1592], lumberyards[1592]}), .bottom({trees[1593], lumberyards[1593]}), .bottom_right({trees[1594], lumberyards[1594]}), .init(2'b00), .state({trees[1543], lumberyards[1543]}));
acre acre_30_44 (.clk(clk), .en(en), .top_left({trees[1493], lumberyards[1493]}), .top({trees[1494], lumberyards[1494]}), .top_right({trees[1495], lumberyards[1495]}), .left({trees[1543], lumberyards[1543]}), .right({trees[1545], lumberyards[1545]}), .bottom_left({trees[1593], lumberyards[1593]}), .bottom({trees[1594], lumberyards[1594]}), .bottom_right({trees[1595], lumberyards[1595]}), .init(2'b00), .state({trees[1544], lumberyards[1544]}));
acre acre_30_45 (.clk(clk), .en(en), .top_left({trees[1494], lumberyards[1494]}), .top({trees[1495], lumberyards[1495]}), .top_right({trees[1496], lumberyards[1496]}), .left({trees[1544], lumberyards[1544]}), .right({trees[1546], lumberyards[1546]}), .bottom_left({trees[1594], lumberyards[1594]}), .bottom({trees[1595], lumberyards[1595]}), .bottom_right({trees[1596], lumberyards[1596]}), .init(2'b00), .state({trees[1545], lumberyards[1545]}));
acre acre_30_46 (.clk(clk), .en(en), .top_left({trees[1495], lumberyards[1495]}), .top({trees[1496], lumberyards[1496]}), .top_right({trees[1497], lumberyards[1497]}), .left({trees[1545], lumberyards[1545]}), .right({trees[1547], lumberyards[1547]}), .bottom_left({trees[1595], lumberyards[1595]}), .bottom({trees[1596], lumberyards[1596]}), .bottom_right({trees[1597], lumberyards[1597]}), .init(2'b10), .state({trees[1546], lumberyards[1546]}));
acre acre_30_47 (.clk(clk), .en(en), .top_left({trees[1496], lumberyards[1496]}), .top({trees[1497], lumberyards[1497]}), .top_right({trees[1498], lumberyards[1498]}), .left({trees[1546], lumberyards[1546]}), .right({trees[1548], lumberyards[1548]}), .bottom_left({trees[1596], lumberyards[1596]}), .bottom({trees[1597], lumberyards[1597]}), .bottom_right({trees[1598], lumberyards[1598]}), .init(2'b00), .state({trees[1547], lumberyards[1547]}));
acre acre_30_48 (.clk(clk), .en(en), .top_left({trees[1497], lumberyards[1497]}), .top({trees[1498], lumberyards[1498]}), .top_right({trees[1499], lumberyards[1499]}), .left({trees[1547], lumberyards[1547]}), .right({trees[1549], lumberyards[1549]}), .bottom_left({trees[1597], lumberyards[1597]}), .bottom({trees[1598], lumberyards[1598]}), .bottom_right({trees[1599], lumberyards[1599]}), .init(2'b00), .state({trees[1548], lumberyards[1548]}));
acre acre_30_49 (.clk(clk), .en(en), .top_left({trees[1498], lumberyards[1498]}), .top({trees[1499], lumberyards[1499]}), .top_right(2'b0), .left({trees[1548], lumberyards[1548]}), .right(2'b0), .bottom_left({trees[1598], lumberyards[1598]}), .bottom({trees[1599], lumberyards[1599]}), .bottom_right(2'b0), .init(2'b01), .state({trees[1549], lumberyards[1549]}));
acre acre_31_0 (.clk(clk), .en(en), .top_left(2'b0), .top({trees[1500], lumberyards[1500]}), .top_right({trees[1501], lumberyards[1501]}), .left(2'b0), .right({trees[1551], lumberyards[1551]}), .bottom_left(2'b0), .bottom({trees[1600], lumberyards[1600]}), .bottom_right({trees[1601], lumberyards[1601]}), .init(2'b10), .state({trees[1550], lumberyards[1550]}));
acre acre_31_1 (.clk(clk), .en(en), .top_left({trees[1500], lumberyards[1500]}), .top({trees[1501], lumberyards[1501]}), .top_right({trees[1502], lumberyards[1502]}), .left({trees[1550], lumberyards[1550]}), .right({trees[1552], lumberyards[1552]}), .bottom_left({trees[1600], lumberyards[1600]}), .bottom({trees[1601], lumberyards[1601]}), .bottom_right({trees[1602], lumberyards[1602]}), .init(2'b00), .state({trees[1551], lumberyards[1551]}));
acre acre_31_2 (.clk(clk), .en(en), .top_left({trees[1501], lumberyards[1501]}), .top({trees[1502], lumberyards[1502]}), .top_right({trees[1503], lumberyards[1503]}), .left({trees[1551], lumberyards[1551]}), .right({trees[1553], lumberyards[1553]}), .bottom_left({trees[1601], lumberyards[1601]}), .bottom({trees[1602], lumberyards[1602]}), .bottom_right({trees[1603], lumberyards[1603]}), .init(2'b00), .state({trees[1552], lumberyards[1552]}));
acre acre_31_3 (.clk(clk), .en(en), .top_left({trees[1502], lumberyards[1502]}), .top({trees[1503], lumberyards[1503]}), .top_right({trees[1504], lumberyards[1504]}), .left({trees[1552], lumberyards[1552]}), .right({trees[1554], lumberyards[1554]}), .bottom_left({trees[1602], lumberyards[1602]}), .bottom({trees[1603], lumberyards[1603]}), .bottom_right({trees[1604], lumberyards[1604]}), .init(2'b00), .state({trees[1553], lumberyards[1553]}));
acre acre_31_4 (.clk(clk), .en(en), .top_left({trees[1503], lumberyards[1503]}), .top({trees[1504], lumberyards[1504]}), .top_right({trees[1505], lumberyards[1505]}), .left({trees[1553], lumberyards[1553]}), .right({trees[1555], lumberyards[1555]}), .bottom_left({trees[1603], lumberyards[1603]}), .bottom({trees[1604], lumberyards[1604]}), .bottom_right({trees[1605], lumberyards[1605]}), .init(2'b00), .state({trees[1554], lumberyards[1554]}));
acre acre_31_5 (.clk(clk), .en(en), .top_left({trees[1504], lumberyards[1504]}), .top({trees[1505], lumberyards[1505]}), .top_right({trees[1506], lumberyards[1506]}), .left({trees[1554], lumberyards[1554]}), .right({trees[1556], lumberyards[1556]}), .bottom_left({trees[1604], lumberyards[1604]}), .bottom({trees[1605], lumberyards[1605]}), .bottom_right({trees[1606], lumberyards[1606]}), .init(2'b00), .state({trees[1555], lumberyards[1555]}));
acre acre_31_6 (.clk(clk), .en(en), .top_left({trees[1505], lumberyards[1505]}), .top({trees[1506], lumberyards[1506]}), .top_right({trees[1507], lumberyards[1507]}), .left({trees[1555], lumberyards[1555]}), .right({trees[1557], lumberyards[1557]}), .bottom_left({trees[1605], lumberyards[1605]}), .bottom({trees[1606], lumberyards[1606]}), .bottom_right({trees[1607], lumberyards[1607]}), .init(2'b00), .state({trees[1556], lumberyards[1556]}));
acre acre_31_7 (.clk(clk), .en(en), .top_left({trees[1506], lumberyards[1506]}), .top({trees[1507], lumberyards[1507]}), .top_right({trees[1508], lumberyards[1508]}), .left({trees[1556], lumberyards[1556]}), .right({trees[1558], lumberyards[1558]}), .bottom_left({trees[1606], lumberyards[1606]}), .bottom({trees[1607], lumberyards[1607]}), .bottom_right({trees[1608], lumberyards[1608]}), .init(2'b00), .state({trees[1557], lumberyards[1557]}));
acre acre_31_8 (.clk(clk), .en(en), .top_left({trees[1507], lumberyards[1507]}), .top({trees[1508], lumberyards[1508]}), .top_right({trees[1509], lumberyards[1509]}), .left({trees[1557], lumberyards[1557]}), .right({trees[1559], lumberyards[1559]}), .bottom_left({trees[1607], lumberyards[1607]}), .bottom({trees[1608], lumberyards[1608]}), .bottom_right({trees[1609], lumberyards[1609]}), .init(2'b00), .state({trees[1558], lumberyards[1558]}));
acre acre_31_9 (.clk(clk), .en(en), .top_left({trees[1508], lumberyards[1508]}), .top({trees[1509], lumberyards[1509]}), .top_right({trees[1510], lumberyards[1510]}), .left({trees[1558], lumberyards[1558]}), .right({trees[1560], lumberyards[1560]}), .bottom_left({trees[1608], lumberyards[1608]}), .bottom({trees[1609], lumberyards[1609]}), .bottom_right({trees[1610], lumberyards[1610]}), .init(2'b00), .state({trees[1559], lumberyards[1559]}));
acre acre_31_10 (.clk(clk), .en(en), .top_left({trees[1509], lumberyards[1509]}), .top({trees[1510], lumberyards[1510]}), .top_right({trees[1511], lumberyards[1511]}), .left({trees[1559], lumberyards[1559]}), .right({trees[1561], lumberyards[1561]}), .bottom_left({trees[1609], lumberyards[1609]}), .bottom({trees[1610], lumberyards[1610]}), .bottom_right({trees[1611], lumberyards[1611]}), .init(2'b01), .state({trees[1560], lumberyards[1560]}));
acre acre_31_11 (.clk(clk), .en(en), .top_left({trees[1510], lumberyards[1510]}), .top({trees[1511], lumberyards[1511]}), .top_right({trees[1512], lumberyards[1512]}), .left({trees[1560], lumberyards[1560]}), .right({trees[1562], lumberyards[1562]}), .bottom_left({trees[1610], lumberyards[1610]}), .bottom({trees[1611], lumberyards[1611]}), .bottom_right({trees[1612], lumberyards[1612]}), .init(2'b00), .state({trees[1561], lumberyards[1561]}));
acre acre_31_12 (.clk(clk), .en(en), .top_left({trees[1511], lumberyards[1511]}), .top({trees[1512], lumberyards[1512]}), .top_right({trees[1513], lumberyards[1513]}), .left({trees[1561], lumberyards[1561]}), .right({trees[1563], lumberyards[1563]}), .bottom_left({trees[1611], lumberyards[1611]}), .bottom({trees[1612], lumberyards[1612]}), .bottom_right({trees[1613], lumberyards[1613]}), .init(2'b10), .state({trees[1562], lumberyards[1562]}));
acre acre_31_13 (.clk(clk), .en(en), .top_left({trees[1512], lumberyards[1512]}), .top({trees[1513], lumberyards[1513]}), .top_right({trees[1514], lumberyards[1514]}), .left({trees[1562], lumberyards[1562]}), .right({trees[1564], lumberyards[1564]}), .bottom_left({trees[1612], lumberyards[1612]}), .bottom({trees[1613], lumberyards[1613]}), .bottom_right({trees[1614], lumberyards[1614]}), .init(2'b10), .state({trees[1563], lumberyards[1563]}));
acre acre_31_14 (.clk(clk), .en(en), .top_left({trees[1513], lumberyards[1513]}), .top({trees[1514], lumberyards[1514]}), .top_right({trees[1515], lumberyards[1515]}), .left({trees[1563], lumberyards[1563]}), .right({trees[1565], lumberyards[1565]}), .bottom_left({trees[1613], lumberyards[1613]}), .bottom({trees[1614], lumberyards[1614]}), .bottom_right({trees[1615], lumberyards[1615]}), .init(2'b00), .state({trees[1564], lumberyards[1564]}));
acre acre_31_15 (.clk(clk), .en(en), .top_left({trees[1514], lumberyards[1514]}), .top({trees[1515], lumberyards[1515]}), .top_right({trees[1516], lumberyards[1516]}), .left({trees[1564], lumberyards[1564]}), .right({trees[1566], lumberyards[1566]}), .bottom_left({trees[1614], lumberyards[1614]}), .bottom({trees[1615], lumberyards[1615]}), .bottom_right({trees[1616], lumberyards[1616]}), .init(2'b00), .state({trees[1565], lumberyards[1565]}));
acre acre_31_16 (.clk(clk), .en(en), .top_left({trees[1515], lumberyards[1515]}), .top({trees[1516], lumberyards[1516]}), .top_right({trees[1517], lumberyards[1517]}), .left({trees[1565], lumberyards[1565]}), .right({trees[1567], lumberyards[1567]}), .bottom_left({trees[1615], lumberyards[1615]}), .bottom({trees[1616], lumberyards[1616]}), .bottom_right({trees[1617], lumberyards[1617]}), .init(2'b00), .state({trees[1566], lumberyards[1566]}));
acre acre_31_17 (.clk(clk), .en(en), .top_left({trees[1516], lumberyards[1516]}), .top({trees[1517], lumberyards[1517]}), .top_right({trees[1518], lumberyards[1518]}), .left({trees[1566], lumberyards[1566]}), .right({trees[1568], lumberyards[1568]}), .bottom_left({trees[1616], lumberyards[1616]}), .bottom({trees[1617], lumberyards[1617]}), .bottom_right({trees[1618], lumberyards[1618]}), .init(2'b00), .state({trees[1567], lumberyards[1567]}));
acre acre_31_18 (.clk(clk), .en(en), .top_left({trees[1517], lumberyards[1517]}), .top({trees[1518], lumberyards[1518]}), .top_right({trees[1519], lumberyards[1519]}), .left({trees[1567], lumberyards[1567]}), .right({trees[1569], lumberyards[1569]}), .bottom_left({trees[1617], lumberyards[1617]}), .bottom({trees[1618], lumberyards[1618]}), .bottom_right({trees[1619], lumberyards[1619]}), .init(2'b00), .state({trees[1568], lumberyards[1568]}));
acre acre_31_19 (.clk(clk), .en(en), .top_left({trees[1518], lumberyards[1518]}), .top({trees[1519], lumberyards[1519]}), .top_right({trees[1520], lumberyards[1520]}), .left({trees[1568], lumberyards[1568]}), .right({trees[1570], lumberyards[1570]}), .bottom_left({trees[1618], lumberyards[1618]}), .bottom({trees[1619], lumberyards[1619]}), .bottom_right({trees[1620], lumberyards[1620]}), .init(2'b01), .state({trees[1569], lumberyards[1569]}));
acre acre_31_20 (.clk(clk), .en(en), .top_left({trees[1519], lumberyards[1519]}), .top({trees[1520], lumberyards[1520]}), .top_right({trees[1521], lumberyards[1521]}), .left({trees[1569], lumberyards[1569]}), .right({trees[1571], lumberyards[1571]}), .bottom_left({trees[1619], lumberyards[1619]}), .bottom({trees[1620], lumberyards[1620]}), .bottom_right({trees[1621], lumberyards[1621]}), .init(2'b00), .state({trees[1570], lumberyards[1570]}));
acre acre_31_21 (.clk(clk), .en(en), .top_left({trees[1520], lumberyards[1520]}), .top({trees[1521], lumberyards[1521]}), .top_right({trees[1522], lumberyards[1522]}), .left({trees[1570], lumberyards[1570]}), .right({trees[1572], lumberyards[1572]}), .bottom_left({trees[1620], lumberyards[1620]}), .bottom({trees[1621], lumberyards[1621]}), .bottom_right({trees[1622], lumberyards[1622]}), .init(2'b00), .state({trees[1571], lumberyards[1571]}));
acre acre_31_22 (.clk(clk), .en(en), .top_left({trees[1521], lumberyards[1521]}), .top({trees[1522], lumberyards[1522]}), .top_right({trees[1523], lumberyards[1523]}), .left({trees[1571], lumberyards[1571]}), .right({trees[1573], lumberyards[1573]}), .bottom_left({trees[1621], lumberyards[1621]}), .bottom({trees[1622], lumberyards[1622]}), .bottom_right({trees[1623], lumberyards[1623]}), .init(2'b00), .state({trees[1572], lumberyards[1572]}));
acre acre_31_23 (.clk(clk), .en(en), .top_left({trees[1522], lumberyards[1522]}), .top({trees[1523], lumberyards[1523]}), .top_right({trees[1524], lumberyards[1524]}), .left({trees[1572], lumberyards[1572]}), .right({trees[1574], lumberyards[1574]}), .bottom_left({trees[1622], lumberyards[1622]}), .bottom({trees[1623], lumberyards[1623]}), .bottom_right({trees[1624], lumberyards[1624]}), .init(2'b00), .state({trees[1573], lumberyards[1573]}));
acre acre_31_24 (.clk(clk), .en(en), .top_left({trees[1523], lumberyards[1523]}), .top({trees[1524], lumberyards[1524]}), .top_right({trees[1525], lumberyards[1525]}), .left({trees[1573], lumberyards[1573]}), .right({trees[1575], lumberyards[1575]}), .bottom_left({trees[1623], lumberyards[1623]}), .bottom({trees[1624], lumberyards[1624]}), .bottom_right({trees[1625], lumberyards[1625]}), .init(2'b00), .state({trees[1574], lumberyards[1574]}));
acre acre_31_25 (.clk(clk), .en(en), .top_left({trees[1524], lumberyards[1524]}), .top({trees[1525], lumberyards[1525]}), .top_right({trees[1526], lumberyards[1526]}), .left({trees[1574], lumberyards[1574]}), .right({trees[1576], lumberyards[1576]}), .bottom_left({trees[1624], lumberyards[1624]}), .bottom({trees[1625], lumberyards[1625]}), .bottom_right({trees[1626], lumberyards[1626]}), .init(2'b00), .state({trees[1575], lumberyards[1575]}));
acre acre_31_26 (.clk(clk), .en(en), .top_left({trees[1525], lumberyards[1525]}), .top({trees[1526], lumberyards[1526]}), .top_right({trees[1527], lumberyards[1527]}), .left({trees[1575], lumberyards[1575]}), .right({trees[1577], lumberyards[1577]}), .bottom_left({trees[1625], lumberyards[1625]}), .bottom({trees[1626], lumberyards[1626]}), .bottom_right({trees[1627], lumberyards[1627]}), .init(2'b01), .state({trees[1576], lumberyards[1576]}));
acre acre_31_27 (.clk(clk), .en(en), .top_left({trees[1526], lumberyards[1526]}), .top({trees[1527], lumberyards[1527]}), .top_right({trees[1528], lumberyards[1528]}), .left({trees[1576], lumberyards[1576]}), .right({trees[1578], lumberyards[1578]}), .bottom_left({trees[1626], lumberyards[1626]}), .bottom({trees[1627], lumberyards[1627]}), .bottom_right({trees[1628], lumberyards[1628]}), .init(2'b10), .state({trees[1577], lumberyards[1577]}));
acre acre_31_28 (.clk(clk), .en(en), .top_left({trees[1527], lumberyards[1527]}), .top({trees[1528], lumberyards[1528]}), .top_right({trees[1529], lumberyards[1529]}), .left({trees[1577], lumberyards[1577]}), .right({trees[1579], lumberyards[1579]}), .bottom_left({trees[1627], lumberyards[1627]}), .bottom({trees[1628], lumberyards[1628]}), .bottom_right({trees[1629], lumberyards[1629]}), .init(2'b00), .state({trees[1578], lumberyards[1578]}));
acre acre_31_29 (.clk(clk), .en(en), .top_left({trees[1528], lumberyards[1528]}), .top({trees[1529], lumberyards[1529]}), .top_right({trees[1530], lumberyards[1530]}), .left({trees[1578], lumberyards[1578]}), .right({trees[1580], lumberyards[1580]}), .bottom_left({trees[1628], lumberyards[1628]}), .bottom({trees[1629], lumberyards[1629]}), .bottom_right({trees[1630], lumberyards[1630]}), .init(2'b00), .state({trees[1579], lumberyards[1579]}));
acre acre_31_30 (.clk(clk), .en(en), .top_left({trees[1529], lumberyards[1529]}), .top({trees[1530], lumberyards[1530]}), .top_right({trees[1531], lumberyards[1531]}), .left({trees[1579], lumberyards[1579]}), .right({trees[1581], lumberyards[1581]}), .bottom_left({trees[1629], lumberyards[1629]}), .bottom({trees[1630], lumberyards[1630]}), .bottom_right({trees[1631], lumberyards[1631]}), .init(2'b10), .state({trees[1580], lumberyards[1580]}));
acre acre_31_31 (.clk(clk), .en(en), .top_left({trees[1530], lumberyards[1530]}), .top({trees[1531], lumberyards[1531]}), .top_right({trees[1532], lumberyards[1532]}), .left({trees[1580], lumberyards[1580]}), .right({trees[1582], lumberyards[1582]}), .bottom_left({trees[1630], lumberyards[1630]}), .bottom({trees[1631], lumberyards[1631]}), .bottom_right({trees[1632], lumberyards[1632]}), .init(2'b10), .state({trees[1581], lumberyards[1581]}));
acre acre_31_32 (.clk(clk), .en(en), .top_left({trees[1531], lumberyards[1531]}), .top({trees[1532], lumberyards[1532]}), .top_right({trees[1533], lumberyards[1533]}), .left({trees[1581], lumberyards[1581]}), .right({trees[1583], lumberyards[1583]}), .bottom_left({trees[1631], lumberyards[1631]}), .bottom({trees[1632], lumberyards[1632]}), .bottom_right({trees[1633], lumberyards[1633]}), .init(2'b10), .state({trees[1582], lumberyards[1582]}));
acre acre_31_33 (.clk(clk), .en(en), .top_left({trees[1532], lumberyards[1532]}), .top({trees[1533], lumberyards[1533]}), .top_right({trees[1534], lumberyards[1534]}), .left({trees[1582], lumberyards[1582]}), .right({trees[1584], lumberyards[1584]}), .bottom_left({trees[1632], lumberyards[1632]}), .bottom({trees[1633], lumberyards[1633]}), .bottom_right({trees[1634], lumberyards[1634]}), .init(2'b00), .state({trees[1583], lumberyards[1583]}));
acre acre_31_34 (.clk(clk), .en(en), .top_left({trees[1533], lumberyards[1533]}), .top({trees[1534], lumberyards[1534]}), .top_right({trees[1535], lumberyards[1535]}), .left({trees[1583], lumberyards[1583]}), .right({trees[1585], lumberyards[1585]}), .bottom_left({trees[1633], lumberyards[1633]}), .bottom({trees[1634], lumberyards[1634]}), .bottom_right({trees[1635], lumberyards[1635]}), .init(2'b00), .state({trees[1584], lumberyards[1584]}));
acre acre_31_35 (.clk(clk), .en(en), .top_left({trees[1534], lumberyards[1534]}), .top({trees[1535], lumberyards[1535]}), .top_right({trees[1536], lumberyards[1536]}), .left({trees[1584], lumberyards[1584]}), .right({trees[1586], lumberyards[1586]}), .bottom_left({trees[1634], lumberyards[1634]}), .bottom({trees[1635], lumberyards[1635]}), .bottom_right({trees[1636], lumberyards[1636]}), .init(2'b00), .state({trees[1585], lumberyards[1585]}));
acre acre_31_36 (.clk(clk), .en(en), .top_left({trees[1535], lumberyards[1535]}), .top({trees[1536], lumberyards[1536]}), .top_right({trees[1537], lumberyards[1537]}), .left({trees[1585], lumberyards[1585]}), .right({trees[1587], lumberyards[1587]}), .bottom_left({trees[1635], lumberyards[1635]}), .bottom({trees[1636], lumberyards[1636]}), .bottom_right({trees[1637], lumberyards[1637]}), .init(2'b00), .state({trees[1586], lumberyards[1586]}));
acre acre_31_37 (.clk(clk), .en(en), .top_left({trees[1536], lumberyards[1536]}), .top({trees[1537], lumberyards[1537]}), .top_right({trees[1538], lumberyards[1538]}), .left({trees[1586], lumberyards[1586]}), .right({trees[1588], lumberyards[1588]}), .bottom_left({trees[1636], lumberyards[1636]}), .bottom({trees[1637], lumberyards[1637]}), .bottom_right({trees[1638], lumberyards[1638]}), .init(2'b00), .state({trees[1587], lumberyards[1587]}));
acre acre_31_38 (.clk(clk), .en(en), .top_left({trees[1537], lumberyards[1537]}), .top({trees[1538], lumberyards[1538]}), .top_right({trees[1539], lumberyards[1539]}), .left({trees[1587], lumberyards[1587]}), .right({trees[1589], lumberyards[1589]}), .bottom_left({trees[1637], lumberyards[1637]}), .bottom({trees[1638], lumberyards[1638]}), .bottom_right({trees[1639], lumberyards[1639]}), .init(2'b00), .state({trees[1588], lumberyards[1588]}));
acre acre_31_39 (.clk(clk), .en(en), .top_left({trees[1538], lumberyards[1538]}), .top({trees[1539], lumberyards[1539]}), .top_right({trees[1540], lumberyards[1540]}), .left({trees[1588], lumberyards[1588]}), .right({trees[1590], lumberyards[1590]}), .bottom_left({trees[1638], lumberyards[1638]}), .bottom({trees[1639], lumberyards[1639]}), .bottom_right({trees[1640], lumberyards[1640]}), .init(2'b01), .state({trees[1589], lumberyards[1589]}));
acre acre_31_40 (.clk(clk), .en(en), .top_left({trees[1539], lumberyards[1539]}), .top({trees[1540], lumberyards[1540]}), .top_right({trees[1541], lumberyards[1541]}), .left({trees[1589], lumberyards[1589]}), .right({trees[1591], lumberyards[1591]}), .bottom_left({trees[1639], lumberyards[1639]}), .bottom({trees[1640], lumberyards[1640]}), .bottom_right({trees[1641], lumberyards[1641]}), .init(2'b01), .state({trees[1590], lumberyards[1590]}));
acre acre_31_41 (.clk(clk), .en(en), .top_left({trees[1540], lumberyards[1540]}), .top({trees[1541], lumberyards[1541]}), .top_right({trees[1542], lumberyards[1542]}), .left({trees[1590], lumberyards[1590]}), .right({trees[1592], lumberyards[1592]}), .bottom_left({trees[1640], lumberyards[1640]}), .bottom({trees[1641], lumberyards[1641]}), .bottom_right({trees[1642], lumberyards[1642]}), .init(2'b00), .state({trees[1591], lumberyards[1591]}));
acre acre_31_42 (.clk(clk), .en(en), .top_left({trees[1541], lumberyards[1541]}), .top({trees[1542], lumberyards[1542]}), .top_right({trees[1543], lumberyards[1543]}), .left({trees[1591], lumberyards[1591]}), .right({trees[1593], lumberyards[1593]}), .bottom_left({trees[1641], lumberyards[1641]}), .bottom({trees[1642], lumberyards[1642]}), .bottom_right({trees[1643], lumberyards[1643]}), .init(2'b00), .state({trees[1592], lumberyards[1592]}));
acre acre_31_43 (.clk(clk), .en(en), .top_left({trees[1542], lumberyards[1542]}), .top({trees[1543], lumberyards[1543]}), .top_right({trees[1544], lumberyards[1544]}), .left({trees[1592], lumberyards[1592]}), .right({trees[1594], lumberyards[1594]}), .bottom_left({trees[1642], lumberyards[1642]}), .bottom({trees[1643], lumberyards[1643]}), .bottom_right({trees[1644], lumberyards[1644]}), .init(2'b00), .state({trees[1593], lumberyards[1593]}));
acre acre_31_44 (.clk(clk), .en(en), .top_left({trees[1543], lumberyards[1543]}), .top({trees[1544], lumberyards[1544]}), .top_right({trees[1545], lumberyards[1545]}), .left({trees[1593], lumberyards[1593]}), .right({trees[1595], lumberyards[1595]}), .bottom_left({trees[1643], lumberyards[1643]}), .bottom({trees[1644], lumberyards[1644]}), .bottom_right({trees[1645], lumberyards[1645]}), .init(2'b10), .state({trees[1594], lumberyards[1594]}));
acre acre_31_45 (.clk(clk), .en(en), .top_left({trees[1544], lumberyards[1544]}), .top({trees[1545], lumberyards[1545]}), .top_right({trees[1546], lumberyards[1546]}), .left({trees[1594], lumberyards[1594]}), .right({trees[1596], lumberyards[1596]}), .bottom_left({trees[1644], lumberyards[1644]}), .bottom({trees[1645], lumberyards[1645]}), .bottom_right({trees[1646], lumberyards[1646]}), .init(2'b01), .state({trees[1595], lumberyards[1595]}));
acre acre_31_46 (.clk(clk), .en(en), .top_left({trees[1545], lumberyards[1545]}), .top({trees[1546], lumberyards[1546]}), .top_right({trees[1547], lumberyards[1547]}), .left({trees[1595], lumberyards[1595]}), .right({trees[1597], lumberyards[1597]}), .bottom_left({trees[1645], lumberyards[1645]}), .bottom({trees[1646], lumberyards[1646]}), .bottom_right({trees[1647], lumberyards[1647]}), .init(2'b10), .state({trees[1596], lumberyards[1596]}));
acre acre_31_47 (.clk(clk), .en(en), .top_left({trees[1546], lumberyards[1546]}), .top({trees[1547], lumberyards[1547]}), .top_right({trees[1548], lumberyards[1548]}), .left({trees[1596], lumberyards[1596]}), .right({trees[1598], lumberyards[1598]}), .bottom_left({trees[1646], lumberyards[1646]}), .bottom({trees[1647], lumberyards[1647]}), .bottom_right({trees[1648], lumberyards[1648]}), .init(2'b00), .state({trees[1597], lumberyards[1597]}));
acre acre_31_48 (.clk(clk), .en(en), .top_left({trees[1547], lumberyards[1547]}), .top({trees[1548], lumberyards[1548]}), .top_right({trees[1549], lumberyards[1549]}), .left({trees[1597], lumberyards[1597]}), .right({trees[1599], lumberyards[1599]}), .bottom_left({trees[1647], lumberyards[1647]}), .bottom({trees[1648], lumberyards[1648]}), .bottom_right({trees[1649], lumberyards[1649]}), .init(2'b00), .state({trees[1598], lumberyards[1598]}));
acre acre_31_49 (.clk(clk), .en(en), .top_left({trees[1548], lumberyards[1548]}), .top({trees[1549], lumberyards[1549]}), .top_right(2'b0), .left({trees[1598], lumberyards[1598]}), .right(2'b0), .bottom_left({trees[1648], lumberyards[1648]}), .bottom({trees[1649], lumberyards[1649]}), .bottom_right(2'b0), .init(2'b00), .state({trees[1599], lumberyards[1599]}));
acre acre_32_0 (.clk(clk), .en(en), .top_left(2'b0), .top({trees[1550], lumberyards[1550]}), .top_right({trees[1551], lumberyards[1551]}), .left(2'b0), .right({trees[1601], lumberyards[1601]}), .bottom_left(2'b0), .bottom({trees[1650], lumberyards[1650]}), .bottom_right({trees[1651], lumberyards[1651]}), .init(2'b00), .state({trees[1600], lumberyards[1600]}));
acre acre_32_1 (.clk(clk), .en(en), .top_left({trees[1550], lumberyards[1550]}), .top({trees[1551], lumberyards[1551]}), .top_right({trees[1552], lumberyards[1552]}), .left({trees[1600], lumberyards[1600]}), .right({trees[1602], lumberyards[1602]}), .bottom_left({trees[1650], lumberyards[1650]}), .bottom({trees[1651], lumberyards[1651]}), .bottom_right({trees[1652], lumberyards[1652]}), .init(2'b10), .state({trees[1601], lumberyards[1601]}));
acre acre_32_2 (.clk(clk), .en(en), .top_left({trees[1551], lumberyards[1551]}), .top({trees[1552], lumberyards[1552]}), .top_right({trees[1553], lumberyards[1553]}), .left({trees[1601], lumberyards[1601]}), .right({trees[1603], lumberyards[1603]}), .bottom_left({trees[1651], lumberyards[1651]}), .bottom({trees[1652], lumberyards[1652]}), .bottom_right({trees[1653], lumberyards[1653]}), .init(2'b00), .state({trees[1602], lumberyards[1602]}));
acre acre_32_3 (.clk(clk), .en(en), .top_left({trees[1552], lumberyards[1552]}), .top({trees[1553], lumberyards[1553]}), .top_right({trees[1554], lumberyards[1554]}), .left({trees[1602], lumberyards[1602]}), .right({trees[1604], lumberyards[1604]}), .bottom_left({trees[1652], lumberyards[1652]}), .bottom({trees[1653], lumberyards[1653]}), .bottom_right({trees[1654], lumberyards[1654]}), .init(2'b10), .state({trees[1603], lumberyards[1603]}));
acre acre_32_4 (.clk(clk), .en(en), .top_left({trees[1553], lumberyards[1553]}), .top({trees[1554], lumberyards[1554]}), .top_right({trees[1555], lumberyards[1555]}), .left({trees[1603], lumberyards[1603]}), .right({trees[1605], lumberyards[1605]}), .bottom_left({trees[1653], lumberyards[1653]}), .bottom({trees[1654], lumberyards[1654]}), .bottom_right({trees[1655], lumberyards[1655]}), .init(2'b10), .state({trees[1604], lumberyards[1604]}));
acre acre_32_5 (.clk(clk), .en(en), .top_left({trees[1554], lumberyards[1554]}), .top({trees[1555], lumberyards[1555]}), .top_right({trees[1556], lumberyards[1556]}), .left({trees[1604], lumberyards[1604]}), .right({trees[1606], lumberyards[1606]}), .bottom_left({trees[1654], lumberyards[1654]}), .bottom({trees[1655], lumberyards[1655]}), .bottom_right({trees[1656], lumberyards[1656]}), .init(2'b00), .state({trees[1605], lumberyards[1605]}));
acre acre_32_6 (.clk(clk), .en(en), .top_left({trees[1555], lumberyards[1555]}), .top({trees[1556], lumberyards[1556]}), .top_right({trees[1557], lumberyards[1557]}), .left({trees[1605], lumberyards[1605]}), .right({trees[1607], lumberyards[1607]}), .bottom_left({trees[1655], lumberyards[1655]}), .bottom({trees[1656], lumberyards[1656]}), .bottom_right({trees[1657], lumberyards[1657]}), .init(2'b00), .state({trees[1606], lumberyards[1606]}));
acre acre_32_7 (.clk(clk), .en(en), .top_left({trees[1556], lumberyards[1556]}), .top({trees[1557], lumberyards[1557]}), .top_right({trees[1558], lumberyards[1558]}), .left({trees[1606], lumberyards[1606]}), .right({trees[1608], lumberyards[1608]}), .bottom_left({trees[1656], lumberyards[1656]}), .bottom({trees[1657], lumberyards[1657]}), .bottom_right({trees[1658], lumberyards[1658]}), .init(2'b01), .state({trees[1607], lumberyards[1607]}));
acre acre_32_8 (.clk(clk), .en(en), .top_left({trees[1557], lumberyards[1557]}), .top({trees[1558], lumberyards[1558]}), .top_right({trees[1559], lumberyards[1559]}), .left({trees[1607], lumberyards[1607]}), .right({trees[1609], lumberyards[1609]}), .bottom_left({trees[1657], lumberyards[1657]}), .bottom({trees[1658], lumberyards[1658]}), .bottom_right({trees[1659], lumberyards[1659]}), .init(2'b00), .state({trees[1608], lumberyards[1608]}));
acre acre_32_9 (.clk(clk), .en(en), .top_left({trees[1558], lumberyards[1558]}), .top({trees[1559], lumberyards[1559]}), .top_right({trees[1560], lumberyards[1560]}), .left({trees[1608], lumberyards[1608]}), .right({trees[1610], lumberyards[1610]}), .bottom_left({trees[1658], lumberyards[1658]}), .bottom({trees[1659], lumberyards[1659]}), .bottom_right({trees[1660], lumberyards[1660]}), .init(2'b00), .state({trees[1609], lumberyards[1609]}));
acre acre_32_10 (.clk(clk), .en(en), .top_left({trees[1559], lumberyards[1559]}), .top({trees[1560], lumberyards[1560]}), .top_right({trees[1561], lumberyards[1561]}), .left({trees[1609], lumberyards[1609]}), .right({trees[1611], lumberyards[1611]}), .bottom_left({trees[1659], lumberyards[1659]}), .bottom({trees[1660], lumberyards[1660]}), .bottom_right({trees[1661], lumberyards[1661]}), .init(2'b00), .state({trees[1610], lumberyards[1610]}));
acre acre_32_11 (.clk(clk), .en(en), .top_left({trees[1560], lumberyards[1560]}), .top({trees[1561], lumberyards[1561]}), .top_right({trees[1562], lumberyards[1562]}), .left({trees[1610], lumberyards[1610]}), .right({trees[1612], lumberyards[1612]}), .bottom_left({trees[1660], lumberyards[1660]}), .bottom({trees[1661], lumberyards[1661]}), .bottom_right({trees[1662], lumberyards[1662]}), .init(2'b10), .state({trees[1611], lumberyards[1611]}));
acre acre_32_12 (.clk(clk), .en(en), .top_left({trees[1561], lumberyards[1561]}), .top({trees[1562], lumberyards[1562]}), .top_right({trees[1563], lumberyards[1563]}), .left({trees[1611], lumberyards[1611]}), .right({trees[1613], lumberyards[1613]}), .bottom_left({trees[1661], lumberyards[1661]}), .bottom({trees[1662], lumberyards[1662]}), .bottom_right({trees[1663], lumberyards[1663]}), .init(2'b00), .state({trees[1612], lumberyards[1612]}));
acre acre_32_13 (.clk(clk), .en(en), .top_left({trees[1562], lumberyards[1562]}), .top({trees[1563], lumberyards[1563]}), .top_right({trees[1564], lumberyards[1564]}), .left({trees[1612], lumberyards[1612]}), .right({trees[1614], lumberyards[1614]}), .bottom_left({trees[1662], lumberyards[1662]}), .bottom({trees[1663], lumberyards[1663]}), .bottom_right({trees[1664], lumberyards[1664]}), .init(2'b00), .state({trees[1613], lumberyards[1613]}));
acre acre_32_14 (.clk(clk), .en(en), .top_left({trees[1563], lumberyards[1563]}), .top({trees[1564], lumberyards[1564]}), .top_right({trees[1565], lumberyards[1565]}), .left({trees[1613], lumberyards[1613]}), .right({trees[1615], lumberyards[1615]}), .bottom_left({trees[1663], lumberyards[1663]}), .bottom({trees[1664], lumberyards[1664]}), .bottom_right({trees[1665], lumberyards[1665]}), .init(2'b10), .state({trees[1614], lumberyards[1614]}));
acre acre_32_15 (.clk(clk), .en(en), .top_left({trees[1564], lumberyards[1564]}), .top({trees[1565], lumberyards[1565]}), .top_right({trees[1566], lumberyards[1566]}), .left({trees[1614], lumberyards[1614]}), .right({trees[1616], lumberyards[1616]}), .bottom_left({trees[1664], lumberyards[1664]}), .bottom({trees[1665], lumberyards[1665]}), .bottom_right({trees[1666], lumberyards[1666]}), .init(2'b00), .state({trees[1615], lumberyards[1615]}));
acre acre_32_16 (.clk(clk), .en(en), .top_left({trees[1565], lumberyards[1565]}), .top({trees[1566], lumberyards[1566]}), .top_right({trees[1567], lumberyards[1567]}), .left({trees[1615], lumberyards[1615]}), .right({trees[1617], lumberyards[1617]}), .bottom_left({trees[1665], lumberyards[1665]}), .bottom({trees[1666], lumberyards[1666]}), .bottom_right({trees[1667], lumberyards[1667]}), .init(2'b00), .state({trees[1616], lumberyards[1616]}));
acre acre_32_17 (.clk(clk), .en(en), .top_left({trees[1566], lumberyards[1566]}), .top({trees[1567], lumberyards[1567]}), .top_right({trees[1568], lumberyards[1568]}), .left({trees[1616], lumberyards[1616]}), .right({trees[1618], lumberyards[1618]}), .bottom_left({trees[1666], lumberyards[1666]}), .bottom({trees[1667], lumberyards[1667]}), .bottom_right({trees[1668], lumberyards[1668]}), .init(2'b00), .state({trees[1617], lumberyards[1617]}));
acre acre_32_18 (.clk(clk), .en(en), .top_left({trees[1567], lumberyards[1567]}), .top({trees[1568], lumberyards[1568]}), .top_right({trees[1569], lumberyards[1569]}), .left({trees[1617], lumberyards[1617]}), .right({trees[1619], lumberyards[1619]}), .bottom_left({trees[1667], lumberyards[1667]}), .bottom({trees[1668], lumberyards[1668]}), .bottom_right({trees[1669], lumberyards[1669]}), .init(2'b00), .state({trees[1618], lumberyards[1618]}));
acre acre_32_19 (.clk(clk), .en(en), .top_left({trees[1568], lumberyards[1568]}), .top({trees[1569], lumberyards[1569]}), .top_right({trees[1570], lumberyards[1570]}), .left({trees[1618], lumberyards[1618]}), .right({trees[1620], lumberyards[1620]}), .bottom_left({trees[1668], lumberyards[1668]}), .bottom({trees[1669], lumberyards[1669]}), .bottom_right({trees[1670], lumberyards[1670]}), .init(2'b00), .state({trees[1619], lumberyards[1619]}));
acre acre_32_20 (.clk(clk), .en(en), .top_left({trees[1569], lumberyards[1569]}), .top({trees[1570], lumberyards[1570]}), .top_right({trees[1571], lumberyards[1571]}), .left({trees[1619], lumberyards[1619]}), .right({trees[1621], lumberyards[1621]}), .bottom_left({trees[1669], lumberyards[1669]}), .bottom({trees[1670], lumberyards[1670]}), .bottom_right({trees[1671], lumberyards[1671]}), .init(2'b00), .state({trees[1620], lumberyards[1620]}));
acre acre_32_21 (.clk(clk), .en(en), .top_left({trees[1570], lumberyards[1570]}), .top({trees[1571], lumberyards[1571]}), .top_right({trees[1572], lumberyards[1572]}), .left({trees[1620], lumberyards[1620]}), .right({trees[1622], lumberyards[1622]}), .bottom_left({trees[1670], lumberyards[1670]}), .bottom({trees[1671], lumberyards[1671]}), .bottom_right({trees[1672], lumberyards[1672]}), .init(2'b01), .state({trees[1621], lumberyards[1621]}));
acre acre_32_22 (.clk(clk), .en(en), .top_left({trees[1571], lumberyards[1571]}), .top({trees[1572], lumberyards[1572]}), .top_right({trees[1573], lumberyards[1573]}), .left({trees[1621], lumberyards[1621]}), .right({trees[1623], lumberyards[1623]}), .bottom_left({trees[1671], lumberyards[1671]}), .bottom({trees[1672], lumberyards[1672]}), .bottom_right({trees[1673], lumberyards[1673]}), .init(2'b00), .state({trees[1622], lumberyards[1622]}));
acre acre_32_23 (.clk(clk), .en(en), .top_left({trees[1572], lumberyards[1572]}), .top({trees[1573], lumberyards[1573]}), .top_right({trees[1574], lumberyards[1574]}), .left({trees[1622], lumberyards[1622]}), .right({trees[1624], lumberyards[1624]}), .bottom_left({trees[1672], lumberyards[1672]}), .bottom({trees[1673], lumberyards[1673]}), .bottom_right({trees[1674], lumberyards[1674]}), .init(2'b00), .state({trees[1623], lumberyards[1623]}));
acre acre_32_24 (.clk(clk), .en(en), .top_left({trees[1573], lumberyards[1573]}), .top({trees[1574], lumberyards[1574]}), .top_right({trees[1575], lumberyards[1575]}), .left({trees[1623], lumberyards[1623]}), .right({trees[1625], lumberyards[1625]}), .bottom_left({trees[1673], lumberyards[1673]}), .bottom({trees[1674], lumberyards[1674]}), .bottom_right({trees[1675], lumberyards[1675]}), .init(2'b00), .state({trees[1624], lumberyards[1624]}));
acre acre_32_25 (.clk(clk), .en(en), .top_left({trees[1574], lumberyards[1574]}), .top({trees[1575], lumberyards[1575]}), .top_right({trees[1576], lumberyards[1576]}), .left({trees[1624], lumberyards[1624]}), .right({trees[1626], lumberyards[1626]}), .bottom_left({trees[1674], lumberyards[1674]}), .bottom({trees[1675], lumberyards[1675]}), .bottom_right({trees[1676], lumberyards[1676]}), .init(2'b00), .state({trees[1625], lumberyards[1625]}));
acre acre_32_26 (.clk(clk), .en(en), .top_left({trees[1575], lumberyards[1575]}), .top({trees[1576], lumberyards[1576]}), .top_right({trees[1577], lumberyards[1577]}), .left({trees[1625], lumberyards[1625]}), .right({trees[1627], lumberyards[1627]}), .bottom_left({trees[1675], lumberyards[1675]}), .bottom({trees[1676], lumberyards[1676]}), .bottom_right({trees[1677], lumberyards[1677]}), .init(2'b00), .state({trees[1626], lumberyards[1626]}));
acre acre_32_27 (.clk(clk), .en(en), .top_left({trees[1576], lumberyards[1576]}), .top({trees[1577], lumberyards[1577]}), .top_right({trees[1578], lumberyards[1578]}), .left({trees[1626], lumberyards[1626]}), .right({trees[1628], lumberyards[1628]}), .bottom_left({trees[1676], lumberyards[1676]}), .bottom({trees[1677], lumberyards[1677]}), .bottom_right({trees[1678], lumberyards[1678]}), .init(2'b00), .state({trees[1627], lumberyards[1627]}));
acre acre_32_28 (.clk(clk), .en(en), .top_left({trees[1577], lumberyards[1577]}), .top({trees[1578], lumberyards[1578]}), .top_right({trees[1579], lumberyards[1579]}), .left({trees[1627], lumberyards[1627]}), .right({trees[1629], lumberyards[1629]}), .bottom_left({trees[1677], lumberyards[1677]}), .bottom({trees[1678], lumberyards[1678]}), .bottom_right({trees[1679], lumberyards[1679]}), .init(2'b00), .state({trees[1628], lumberyards[1628]}));
acre acre_32_29 (.clk(clk), .en(en), .top_left({trees[1578], lumberyards[1578]}), .top({trees[1579], lumberyards[1579]}), .top_right({trees[1580], lumberyards[1580]}), .left({trees[1628], lumberyards[1628]}), .right({trees[1630], lumberyards[1630]}), .bottom_left({trees[1678], lumberyards[1678]}), .bottom({trees[1679], lumberyards[1679]}), .bottom_right({trees[1680], lumberyards[1680]}), .init(2'b10), .state({trees[1629], lumberyards[1629]}));
acre acre_32_30 (.clk(clk), .en(en), .top_left({trees[1579], lumberyards[1579]}), .top({trees[1580], lumberyards[1580]}), .top_right({trees[1581], lumberyards[1581]}), .left({trees[1629], lumberyards[1629]}), .right({trees[1631], lumberyards[1631]}), .bottom_left({trees[1679], lumberyards[1679]}), .bottom({trees[1680], lumberyards[1680]}), .bottom_right({trees[1681], lumberyards[1681]}), .init(2'b00), .state({trees[1630], lumberyards[1630]}));
acre acre_32_31 (.clk(clk), .en(en), .top_left({trees[1580], lumberyards[1580]}), .top({trees[1581], lumberyards[1581]}), .top_right({trees[1582], lumberyards[1582]}), .left({trees[1630], lumberyards[1630]}), .right({trees[1632], lumberyards[1632]}), .bottom_left({trees[1680], lumberyards[1680]}), .bottom({trees[1681], lumberyards[1681]}), .bottom_right({trees[1682], lumberyards[1682]}), .init(2'b00), .state({trees[1631], lumberyards[1631]}));
acre acre_32_32 (.clk(clk), .en(en), .top_left({trees[1581], lumberyards[1581]}), .top({trees[1582], lumberyards[1582]}), .top_right({trees[1583], lumberyards[1583]}), .left({trees[1631], lumberyards[1631]}), .right({trees[1633], lumberyards[1633]}), .bottom_left({trees[1681], lumberyards[1681]}), .bottom({trees[1682], lumberyards[1682]}), .bottom_right({trees[1683], lumberyards[1683]}), .init(2'b00), .state({trees[1632], lumberyards[1632]}));
acre acre_32_33 (.clk(clk), .en(en), .top_left({trees[1582], lumberyards[1582]}), .top({trees[1583], lumberyards[1583]}), .top_right({trees[1584], lumberyards[1584]}), .left({trees[1632], lumberyards[1632]}), .right({trees[1634], lumberyards[1634]}), .bottom_left({trees[1682], lumberyards[1682]}), .bottom({trees[1683], lumberyards[1683]}), .bottom_right({trees[1684], lumberyards[1684]}), .init(2'b10), .state({trees[1633], lumberyards[1633]}));
acre acre_32_34 (.clk(clk), .en(en), .top_left({trees[1583], lumberyards[1583]}), .top({trees[1584], lumberyards[1584]}), .top_right({trees[1585], lumberyards[1585]}), .left({trees[1633], lumberyards[1633]}), .right({trees[1635], lumberyards[1635]}), .bottom_left({trees[1683], lumberyards[1683]}), .bottom({trees[1684], lumberyards[1684]}), .bottom_right({trees[1685], lumberyards[1685]}), .init(2'b00), .state({trees[1634], lumberyards[1634]}));
acre acre_32_35 (.clk(clk), .en(en), .top_left({trees[1584], lumberyards[1584]}), .top({trees[1585], lumberyards[1585]}), .top_right({trees[1586], lumberyards[1586]}), .left({trees[1634], lumberyards[1634]}), .right({trees[1636], lumberyards[1636]}), .bottom_left({trees[1684], lumberyards[1684]}), .bottom({trees[1685], lumberyards[1685]}), .bottom_right({trees[1686], lumberyards[1686]}), .init(2'b10), .state({trees[1635], lumberyards[1635]}));
acre acre_32_36 (.clk(clk), .en(en), .top_left({trees[1585], lumberyards[1585]}), .top({trees[1586], lumberyards[1586]}), .top_right({trees[1587], lumberyards[1587]}), .left({trees[1635], lumberyards[1635]}), .right({trees[1637], lumberyards[1637]}), .bottom_left({trees[1685], lumberyards[1685]}), .bottom({trees[1686], lumberyards[1686]}), .bottom_right({trees[1687], lumberyards[1687]}), .init(2'b01), .state({trees[1636], lumberyards[1636]}));
acre acre_32_37 (.clk(clk), .en(en), .top_left({trees[1586], lumberyards[1586]}), .top({trees[1587], lumberyards[1587]}), .top_right({trees[1588], lumberyards[1588]}), .left({trees[1636], lumberyards[1636]}), .right({trees[1638], lumberyards[1638]}), .bottom_left({trees[1686], lumberyards[1686]}), .bottom({trees[1687], lumberyards[1687]}), .bottom_right({trees[1688], lumberyards[1688]}), .init(2'b10), .state({trees[1637], lumberyards[1637]}));
acre acre_32_38 (.clk(clk), .en(en), .top_left({trees[1587], lumberyards[1587]}), .top({trees[1588], lumberyards[1588]}), .top_right({trees[1589], lumberyards[1589]}), .left({trees[1637], lumberyards[1637]}), .right({trees[1639], lumberyards[1639]}), .bottom_left({trees[1687], lumberyards[1687]}), .bottom({trees[1688], lumberyards[1688]}), .bottom_right({trees[1689], lumberyards[1689]}), .init(2'b00), .state({trees[1638], lumberyards[1638]}));
acre acre_32_39 (.clk(clk), .en(en), .top_left({trees[1588], lumberyards[1588]}), .top({trees[1589], lumberyards[1589]}), .top_right({trees[1590], lumberyards[1590]}), .left({trees[1638], lumberyards[1638]}), .right({trees[1640], lumberyards[1640]}), .bottom_left({trees[1688], lumberyards[1688]}), .bottom({trees[1689], lumberyards[1689]}), .bottom_right({trees[1690], lumberyards[1690]}), .init(2'b00), .state({trees[1639], lumberyards[1639]}));
acre acre_32_40 (.clk(clk), .en(en), .top_left({trees[1589], lumberyards[1589]}), .top({trees[1590], lumberyards[1590]}), .top_right({trees[1591], lumberyards[1591]}), .left({trees[1639], lumberyards[1639]}), .right({trees[1641], lumberyards[1641]}), .bottom_left({trees[1689], lumberyards[1689]}), .bottom({trees[1690], lumberyards[1690]}), .bottom_right({trees[1691], lumberyards[1691]}), .init(2'b00), .state({trees[1640], lumberyards[1640]}));
acre acre_32_41 (.clk(clk), .en(en), .top_left({trees[1590], lumberyards[1590]}), .top({trees[1591], lumberyards[1591]}), .top_right({trees[1592], lumberyards[1592]}), .left({trees[1640], lumberyards[1640]}), .right({trees[1642], lumberyards[1642]}), .bottom_left({trees[1690], lumberyards[1690]}), .bottom({trees[1691], lumberyards[1691]}), .bottom_right({trees[1692], lumberyards[1692]}), .init(2'b00), .state({trees[1641], lumberyards[1641]}));
acre acre_32_42 (.clk(clk), .en(en), .top_left({trees[1591], lumberyards[1591]}), .top({trees[1592], lumberyards[1592]}), .top_right({trees[1593], lumberyards[1593]}), .left({trees[1641], lumberyards[1641]}), .right({trees[1643], lumberyards[1643]}), .bottom_left({trees[1691], lumberyards[1691]}), .bottom({trees[1692], lumberyards[1692]}), .bottom_right({trees[1693], lumberyards[1693]}), .init(2'b01), .state({trees[1642], lumberyards[1642]}));
acre acre_32_43 (.clk(clk), .en(en), .top_left({trees[1592], lumberyards[1592]}), .top({trees[1593], lumberyards[1593]}), .top_right({trees[1594], lumberyards[1594]}), .left({trees[1642], lumberyards[1642]}), .right({trees[1644], lumberyards[1644]}), .bottom_left({trees[1692], lumberyards[1692]}), .bottom({trees[1693], lumberyards[1693]}), .bottom_right({trees[1694], lumberyards[1694]}), .init(2'b00), .state({trees[1643], lumberyards[1643]}));
acre acre_32_44 (.clk(clk), .en(en), .top_left({trees[1593], lumberyards[1593]}), .top({trees[1594], lumberyards[1594]}), .top_right({trees[1595], lumberyards[1595]}), .left({trees[1643], lumberyards[1643]}), .right({trees[1645], lumberyards[1645]}), .bottom_left({trees[1693], lumberyards[1693]}), .bottom({trees[1694], lumberyards[1694]}), .bottom_right({trees[1695], lumberyards[1695]}), .init(2'b10), .state({trees[1644], lumberyards[1644]}));
acre acre_32_45 (.clk(clk), .en(en), .top_left({trees[1594], lumberyards[1594]}), .top({trees[1595], lumberyards[1595]}), .top_right({trees[1596], lumberyards[1596]}), .left({trees[1644], lumberyards[1644]}), .right({trees[1646], lumberyards[1646]}), .bottom_left({trees[1694], lumberyards[1694]}), .bottom({trees[1695], lumberyards[1695]}), .bottom_right({trees[1696], lumberyards[1696]}), .init(2'b00), .state({trees[1645], lumberyards[1645]}));
acre acre_32_46 (.clk(clk), .en(en), .top_left({trees[1595], lumberyards[1595]}), .top({trees[1596], lumberyards[1596]}), .top_right({trees[1597], lumberyards[1597]}), .left({trees[1645], lumberyards[1645]}), .right({trees[1647], lumberyards[1647]}), .bottom_left({trees[1695], lumberyards[1695]}), .bottom({trees[1696], lumberyards[1696]}), .bottom_right({trees[1697], lumberyards[1697]}), .init(2'b00), .state({trees[1646], lumberyards[1646]}));
acre acre_32_47 (.clk(clk), .en(en), .top_left({trees[1596], lumberyards[1596]}), .top({trees[1597], lumberyards[1597]}), .top_right({trees[1598], lumberyards[1598]}), .left({trees[1646], lumberyards[1646]}), .right({trees[1648], lumberyards[1648]}), .bottom_left({trees[1696], lumberyards[1696]}), .bottom({trees[1697], lumberyards[1697]}), .bottom_right({trees[1698], lumberyards[1698]}), .init(2'b00), .state({trees[1647], lumberyards[1647]}));
acre acre_32_48 (.clk(clk), .en(en), .top_left({trees[1597], lumberyards[1597]}), .top({trees[1598], lumberyards[1598]}), .top_right({trees[1599], lumberyards[1599]}), .left({trees[1647], lumberyards[1647]}), .right({trees[1649], lumberyards[1649]}), .bottom_left({trees[1697], lumberyards[1697]}), .bottom({trees[1698], lumberyards[1698]}), .bottom_right({trees[1699], lumberyards[1699]}), .init(2'b00), .state({trees[1648], lumberyards[1648]}));
acre acre_32_49 (.clk(clk), .en(en), .top_left({trees[1598], lumberyards[1598]}), .top({trees[1599], lumberyards[1599]}), .top_right(2'b0), .left({trees[1648], lumberyards[1648]}), .right(2'b0), .bottom_left({trees[1698], lumberyards[1698]}), .bottom({trees[1699], lumberyards[1699]}), .bottom_right(2'b0), .init(2'b01), .state({trees[1649], lumberyards[1649]}));
acre acre_33_0 (.clk(clk), .en(en), .top_left(2'b0), .top({trees[1600], lumberyards[1600]}), .top_right({trees[1601], lumberyards[1601]}), .left(2'b0), .right({trees[1651], lumberyards[1651]}), .bottom_left(2'b0), .bottom({trees[1700], lumberyards[1700]}), .bottom_right({trees[1701], lumberyards[1701]}), .init(2'b00), .state({trees[1650], lumberyards[1650]}));
acre acre_33_1 (.clk(clk), .en(en), .top_left({trees[1600], lumberyards[1600]}), .top({trees[1601], lumberyards[1601]}), .top_right({trees[1602], lumberyards[1602]}), .left({trees[1650], lumberyards[1650]}), .right({trees[1652], lumberyards[1652]}), .bottom_left({trees[1700], lumberyards[1700]}), .bottom({trees[1701], lumberyards[1701]}), .bottom_right({trees[1702], lumberyards[1702]}), .init(2'b01), .state({trees[1651], lumberyards[1651]}));
acre acre_33_2 (.clk(clk), .en(en), .top_left({trees[1601], lumberyards[1601]}), .top({trees[1602], lumberyards[1602]}), .top_right({trees[1603], lumberyards[1603]}), .left({trees[1651], lumberyards[1651]}), .right({trees[1653], lumberyards[1653]}), .bottom_left({trees[1701], lumberyards[1701]}), .bottom({trees[1702], lumberyards[1702]}), .bottom_right({trees[1703], lumberyards[1703]}), .init(2'b00), .state({trees[1652], lumberyards[1652]}));
acre acre_33_3 (.clk(clk), .en(en), .top_left({trees[1602], lumberyards[1602]}), .top({trees[1603], lumberyards[1603]}), .top_right({trees[1604], lumberyards[1604]}), .left({trees[1652], lumberyards[1652]}), .right({trees[1654], lumberyards[1654]}), .bottom_left({trees[1702], lumberyards[1702]}), .bottom({trees[1703], lumberyards[1703]}), .bottom_right({trees[1704], lumberyards[1704]}), .init(2'b00), .state({trees[1653], lumberyards[1653]}));
acre acre_33_4 (.clk(clk), .en(en), .top_left({trees[1603], lumberyards[1603]}), .top({trees[1604], lumberyards[1604]}), .top_right({trees[1605], lumberyards[1605]}), .left({trees[1653], lumberyards[1653]}), .right({trees[1655], lumberyards[1655]}), .bottom_left({trees[1703], lumberyards[1703]}), .bottom({trees[1704], lumberyards[1704]}), .bottom_right({trees[1705], lumberyards[1705]}), .init(2'b00), .state({trees[1654], lumberyards[1654]}));
acre acre_33_5 (.clk(clk), .en(en), .top_left({trees[1604], lumberyards[1604]}), .top({trees[1605], lumberyards[1605]}), .top_right({trees[1606], lumberyards[1606]}), .left({trees[1654], lumberyards[1654]}), .right({trees[1656], lumberyards[1656]}), .bottom_left({trees[1704], lumberyards[1704]}), .bottom({trees[1705], lumberyards[1705]}), .bottom_right({trees[1706], lumberyards[1706]}), .init(2'b00), .state({trees[1655], lumberyards[1655]}));
acre acre_33_6 (.clk(clk), .en(en), .top_left({trees[1605], lumberyards[1605]}), .top({trees[1606], lumberyards[1606]}), .top_right({trees[1607], lumberyards[1607]}), .left({trees[1655], lumberyards[1655]}), .right({trees[1657], lumberyards[1657]}), .bottom_left({trees[1705], lumberyards[1705]}), .bottom({trees[1706], lumberyards[1706]}), .bottom_right({trees[1707], lumberyards[1707]}), .init(2'b00), .state({trees[1656], lumberyards[1656]}));
acre acre_33_7 (.clk(clk), .en(en), .top_left({trees[1606], lumberyards[1606]}), .top({trees[1607], lumberyards[1607]}), .top_right({trees[1608], lumberyards[1608]}), .left({trees[1656], lumberyards[1656]}), .right({trees[1658], lumberyards[1658]}), .bottom_left({trees[1706], lumberyards[1706]}), .bottom({trees[1707], lumberyards[1707]}), .bottom_right({trees[1708], lumberyards[1708]}), .init(2'b00), .state({trees[1657], lumberyards[1657]}));
acre acre_33_8 (.clk(clk), .en(en), .top_left({trees[1607], lumberyards[1607]}), .top({trees[1608], lumberyards[1608]}), .top_right({trees[1609], lumberyards[1609]}), .left({trees[1657], lumberyards[1657]}), .right({trees[1659], lumberyards[1659]}), .bottom_left({trees[1707], lumberyards[1707]}), .bottom({trees[1708], lumberyards[1708]}), .bottom_right({trees[1709], lumberyards[1709]}), .init(2'b01), .state({trees[1658], lumberyards[1658]}));
acre acre_33_9 (.clk(clk), .en(en), .top_left({trees[1608], lumberyards[1608]}), .top({trees[1609], lumberyards[1609]}), .top_right({trees[1610], lumberyards[1610]}), .left({trees[1658], lumberyards[1658]}), .right({trees[1660], lumberyards[1660]}), .bottom_left({trees[1708], lumberyards[1708]}), .bottom({trees[1709], lumberyards[1709]}), .bottom_right({trees[1710], lumberyards[1710]}), .init(2'b00), .state({trees[1659], lumberyards[1659]}));
acre acre_33_10 (.clk(clk), .en(en), .top_left({trees[1609], lumberyards[1609]}), .top({trees[1610], lumberyards[1610]}), .top_right({trees[1611], lumberyards[1611]}), .left({trees[1659], lumberyards[1659]}), .right({trees[1661], lumberyards[1661]}), .bottom_left({trees[1709], lumberyards[1709]}), .bottom({trees[1710], lumberyards[1710]}), .bottom_right({trees[1711], lumberyards[1711]}), .init(2'b00), .state({trees[1660], lumberyards[1660]}));
acre acre_33_11 (.clk(clk), .en(en), .top_left({trees[1610], lumberyards[1610]}), .top({trees[1611], lumberyards[1611]}), .top_right({trees[1612], lumberyards[1612]}), .left({trees[1660], lumberyards[1660]}), .right({trees[1662], lumberyards[1662]}), .bottom_left({trees[1710], lumberyards[1710]}), .bottom({trees[1711], lumberyards[1711]}), .bottom_right({trees[1712], lumberyards[1712]}), .init(2'b00), .state({trees[1661], lumberyards[1661]}));
acre acre_33_12 (.clk(clk), .en(en), .top_left({trees[1611], lumberyards[1611]}), .top({trees[1612], lumberyards[1612]}), .top_right({trees[1613], lumberyards[1613]}), .left({trees[1661], lumberyards[1661]}), .right({trees[1663], lumberyards[1663]}), .bottom_left({trees[1711], lumberyards[1711]}), .bottom({trees[1712], lumberyards[1712]}), .bottom_right({trees[1713], lumberyards[1713]}), .init(2'b00), .state({trees[1662], lumberyards[1662]}));
acre acre_33_13 (.clk(clk), .en(en), .top_left({trees[1612], lumberyards[1612]}), .top({trees[1613], lumberyards[1613]}), .top_right({trees[1614], lumberyards[1614]}), .left({trees[1662], lumberyards[1662]}), .right({trees[1664], lumberyards[1664]}), .bottom_left({trees[1712], lumberyards[1712]}), .bottom({trees[1713], lumberyards[1713]}), .bottom_right({trees[1714], lumberyards[1714]}), .init(2'b00), .state({trees[1663], lumberyards[1663]}));
acre acre_33_14 (.clk(clk), .en(en), .top_left({trees[1613], lumberyards[1613]}), .top({trees[1614], lumberyards[1614]}), .top_right({trees[1615], lumberyards[1615]}), .left({trees[1663], lumberyards[1663]}), .right({trees[1665], lumberyards[1665]}), .bottom_left({trees[1713], lumberyards[1713]}), .bottom({trees[1714], lumberyards[1714]}), .bottom_right({trees[1715], lumberyards[1715]}), .init(2'b10), .state({trees[1664], lumberyards[1664]}));
acre acre_33_15 (.clk(clk), .en(en), .top_left({trees[1614], lumberyards[1614]}), .top({trees[1615], lumberyards[1615]}), .top_right({trees[1616], lumberyards[1616]}), .left({trees[1664], lumberyards[1664]}), .right({trees[1666], lumberyards[1666]}), .bottom_left({trees[1714], lumberyards[1714]}), .bottom({trees[1715], lumberyards[1715]}), .bottom_right({trees[1716], lumberyards[1716]}), .init(2'b10), .state({trees[1665], lumberyards[1665]}));
acre acre_33_16 (.clk(clk), .en(en), .top_left({trees[1615], lumberyards[1615]}), .top({trees[1616], lumberyards[1616]}), .top_right({trees[1617], lumberyards[1617]}), .left({trees[1665], lumberyards[1665]}), .right({trees[1667], lumberyards[1667]}), .bottom_left({trees[1715], lumberyards[1715]}), .bottom({trees[1716], lumberyards[1716]}), .bottom_right({trees[1717], lumberyards[1717]}), .init(2'b00), .state({trees[1666], lumberyards[1666]}));
acre acre_33_17 (.clk(clk), .en(en), .top_left({trees[1616], lumberyards[1616]}), .top({trees[1617], lumberyards[1617]}), .top_right({trees[1618], lumberyards[1618]}), .left({trees[1666], lumberyards[1666]}), .right({trees[1668], lumberyards[1668]}), .bottom_left({trees[1716], lumberyards[1716]}), .bottom({trees[1717], lumberyards[1717]}), .bottom_right({trees[1718], lumberyards[1718]}), .init(2'b10), .state({trees[1667], lumberyards[1667]}));
acre acre_33_18 (.clk(clk), .en(en), .top_left({trees[1617], lumberyards[1617]}), .top({trees[1618], lumberyards[1618]}), .top_right({trees[1619], lumberyards[1619]}), .left({trees[1667], lumberyards[1667]}), .right({trees[1669], lumberyards[1669]}), .bottom_left({trees[1717], lumberyards[1717]}), .bottom({trees[1718], lumberyards[1718]}), .bottom_right({trees[1719], lumberyards[1719]}), .init(2'b00), .state({trees[1668], lumberyards[1668]}));
acre acre_33_19 (.clk(clk), .en(en), .top_left({trees[1618], lumberyards[1618]}), .top({trees[1619], lumberyards[1619]}), .top_right({trees[1620], lumberyards[1620]}), .left({trees[1668], lumberyards[1668]}), .right({trees[1670], lumberyards[1670]}), .bottom_left({trees[1718], lumberyards[1718]}), .bottom({trees[1719], lumberyards[1719]}), .bottom_right({trees[1720], lumberyards[1720]}), .init(2'b00), .state({trees[1669], lumberyards[1669]}));
acre acre_33_20 (.clk(clk), .en(en), .top_left({trees[1619], lumberyards[1619]}), .top({trees[1620], lumberyards[1620]}), .top_right({trees[1621], lumberyards[1621]}), .left({trees[1669], lumberyards[1669]}), .right({trees[1671], lumberyards[1671]}), .bottom_left({trees[1719], lumberyards[1719]}), .bottom({trees[1720], lumberyards[1720]}), .bottom_right({trees[1721], lumberyards[1721]}), .init(2'b00), .state({trees[1670], lumberyards[1670]}));
acre acre_33_21 (.clk(clk), .en(en), .top_left({trees[1620], lumberyards[1620]}), .top({trees[1621], lumberyards[1621]}), .top_right({trees[1622], lumberyards[1622]}), .left({trees[1670], lumberyards[1670]}), .right({trees[1672], lumberyards[1672]}), .bottom_left({trees[1720], lumberyards[1720]}), .bottom({trees[1721], lumberyards[1721]}), .bottom_right({trees[1722], lumberyards[1722]}), .init(2'b00), .state({trees[1671], lumberyards[1671]}));
acre acre_33_22 (.clk(clk), .en(en), .top_left({trees[1621], lumberyards[1621]}), .top({trees[1622], lumberyards[1622]}), .top_right({trees[1623], lumberyards[1623]}), .left({trees[1671], lumberyards[1671]}), .right({trees[1673], lumberyards[1673]}), .bottom_left({trees[1721], lumberyards[1721]}), .bottom({trees[1722], lumberyards[1722]}), .bottom_right({trees[1723], lumberyards[1723]}), .init(2'b00), .state({trees[1672], lumberyards[1672]}));
acre acre_33_23 (.clk(clk), .en(en), .top_left({trees[1622], lumberyards[1622]}), .top({trees[1623], lumberyards[1623]}), .top_right({trees[1624], lumberyards[1624]}), .left({trees[1672], lumberyards[1672]}), .right({trees[1674], lumberyards[1674]}), .bottom_left({trees[1722], lumberyards[1722]}), .bottom({trees[1723], lumberyards[1723]}), .bottom_right({trees[1724], lumberyards[1724]}), .init(2'b00), .state({trees[1673], lumberyards[1673]}));
acre acre_33_24 (.clk(clk), .en(en), .top_left({trees[1623], lumberyards[1623]}), .top({trees[1624], lumberyards[1624]}), .top_right({trees[1625], lumberyards[1625]}), .left({trees[1673], lumberyards[1673]}), .right({trees[1675], lumberyards[1675]}), .bottom_left({trees[1723], lumberyards[1723]}), .bottom({trees[1724], lumberyards[1724]}), .bottom_right({trees[1725], lumberyards[1725]}), .init(2'b00), .state({trees[1674], lumberyards[1674]}));
acre acre_33_25 (.clk(clk), .en(en), .top_left({trees[1624], lumberyards[1624]}), .top({trees[1625], lumberyards[1625]}), .top_right({trees[1626], lumberyards[1626]}), .left({trees[1674], lumberyards[1674]}), .right({trees[1676], lumberyards[1676]}), .bottom_left({trees[1724], lumberyards[1724]}), .bottom({trees[1725], lumberyards[1725]}), .bottom_right({trees[1726], lumberyards[1726]}), .init(2'b10), .state({trees[1675], lumberyards[1675]}));
acre acre_33_26 (.clk(clk), .en(en), .top_left({trees[1625], lumberyards[1625]}), .top({trees[1626], lumberyards[1626]}), .top_right({trees[1627], lumberyards[1627]}), .left({trees[1675], lumberyards[1675]}), .right({trees[1677], lumberyards[1677]}), .bottom_left({trees[1725], lumberyards[1725]}), .bottom({trees[1726], lumberyards[1726]}), .bottom_right({trees[1727], lumberyards[1727]}), .init(2'b01), .state({trees[1676], lumberyards[1676]}));
acre acre_33_27 (.clk(clk), .en(en), .top_left({trees[1626], lumberyards[1626]}), .top({trees[1627], lumberyards[1627]}), .top_right({trees[1628], lumberyards[1628]}), .left({trees[1676], lumberyards[1676]}), .right({trees[1678], lumberyards[1678]}), .bottom_left({trees[1726], lumberyards[1726]}), .bottom({trees[1727], lumberyards[1727]}), .bottom_right({trees[1728], lumberyards[1728]}), .init(2'b10), .state({trees[1677], lumberyards[1677]}));
acre acre_33_28 (.clk(clk), .en(en), .top_left({trees[1627], lumberyards[1627]}), .top({trees[1628], lumberyards[1628]}), .top_right({trees[1629], lumberyards[1629]}), .left({trees[1677], lumberyards[1677]}), .right({trees[1679], lumberyards[1679]}), .bottom_left({trees[1727], lumberyards[1727]}), .bottom({trees[1728], lumberyards[1728]}), .bottom_right({trees[1729], lumberyards[1729]}), .init(2'b10), .state({trees[1678], lumberyards[1678]}));
acre acre_33_29 (.clk(clk), .en(en), .top_left({trees[1628], lumberyards[1628]}), .top({trees[1629], lumberyards[1629]}), .top_right({trees[1630], lumberyards[1630]}), .left({trees[1678], lumberyards[1678]}), .right({trees[1680], lumberyards[1680]}), .bottom_left({trees[1728], lumberyards[1728]}), .bottom({trees[1729], lumberyards[1729]}), .bottom_right({trees[1730], lumberyards[1730]}), .init(2'b00), .state({trees[1679], lumberyards[1679]}));
acre acre_33_30 (.clk(clk), .en(en), .top_left({trees[1629], lumberyards[1629]}), .top({trees[1630], lumberyards[1630]}), .top_right({trees[1631], lumberyards[1631]}), .left({trees[1679], lumberyards[1679]}), .right({trees[1681], lumberyards[1681]}), .bottom_left({trees[1729], lumberyards[1729]}), .bottom({trees[1730], lumberyards[1730]}), .bottom_right({trees[1731], lumberyards[1731]}), .init(2'b01), .state({trees[1680], lumberyards[1680]}));
acre acre_33_31 (.clk(clk), .en(en), .top_left({trees[1630], lumberyards[1630]}), .top({trees[1631], lumberyards[1631]}), .top_right({trees[1632], lumberyards[1632]}), .left({trees[1680], lumberyards[1680]}), .right({trees[1682], lumberyards[1682]}), .bottom_left({trees[1730], lumberyards[1730]}), .bottom({trees[1731], lumberyards[1731]}), .bottom_right({trees[1732], lumberyards[1732]}), .init(2'b01), .state({trees[1681], lumberyards[1681]}));
acre acre_33_32 (.clk(clk), .en(en), .top_left({trees[1631], lumberyards[1631]}), .top({trees[1632], lumberyards[1632]}), .top_right({trees[1633], lumberyards[1633]}), .left({trees[1681], lumberyards[1681]}), .right({trees[1683], lumberyards[1683]}), .bottom_left({trees[1731], lumberyards[1731]}), .bottom({trees[1732], lumberyards[1732]}), .bottom_right({trees[1733], lumberyards[1733]}), .init(2'b00), .state({trees[1682], lumberyards[1682]}));
acre acre_33_33 (.clk(clk), .en(en), .top_left({trees[1632], lumberyards[1632]}), .top({trees[1633], lumberyards[1633]}), .top_right({trees[1634], lumberyards[1634]}), .left({trees[1682], lumberyards[1682]}), .right({trees[1684], lumberyards[1684]}), .bottom_left({trees[1732], lumberyards[1732]}), .bottom({trees[1733], lumberyards[1733]}), .bottom_right({trees[1734], lumberyards[1734]}), .init(2'b00), .state({trees[1683], lumberyards[1683]}));
acre acre_33_34 (.clk(clk), .en(en), .top_left({trees[1633], lumberyards[1633]}), .top({trees[1634], lumberyards[1634]}), .top_right({trees[1635], lumberyards[1635]}), .left({trees[1683], lumberyards[1683]}), .right({trees[1685], lumberyards[1685]}), .bottom_left({trees[1733], lumberyards[1733]}), .bottom({trees[1734], lumberyards[1734]}), .bottom_right({trees[1735], lumberyards[1735]}), .init(2'b00), .state({trees[1684], lumberyards[1684]}));
acre acre_33_35 (.clk(clk), .en(en), .top_left({trees[1634], lumberyards[1634]}), .top({trees[1635], lumberyards[1635]}), .top_right({trees[1636], lumberyards[1636]}), .left({trees[1684], lumberyards[1684]}), .right({trees[1686], lumberyards[1686]}), .bottom_left({trees[1734], lumberyards[1734]}), .bottom({trees[1735], lumberyards[1735]}), .bottom_right({trees[1736], lumberyards[1736]}), .init(2'b00), .state({trees[1685], lumberyards[1685]}));
acre acre_33_36 (.clk(clk), .en(en), .top_left({trees[1635], lumberyards[1635]}), .top({trees[1636], lumberyards[1636]}), .top_right({trees[1637], lumberyards[1637]}), .left({trees[1685], lumberyards[1685]}), .right({trees[1687], lumberyards[1687]}), .bottom_left({trees[1735], lumberyards[1735]}), .bottom({trees[1736], lumberyards[1736]}), .bottom_right({trees[1737], lumberyards[1737]}), .init(2'b00), .state({trees[1686], lumberyards[1686]}));
acre acre_33_37 (.clk(clk), .en(en), .top_left({trees[1636], lumberyards[1636]}), .top({trees[1637], lumberyards[1637]}), .top_right({trees[1638], lumberyards[1638]}), .left({trees[1686], lumberyards[1686]}), .right({trees[1688], lumberyards[1688]}), .bottom_left({trees[1736], lumberyards[1736]}), .bottom({trees[1737], lumberyards[1737]}), .bottom_right({trees[1738], lumberyards[1738]}), .init(2'b00), .state({trees[1687], lumberyards[1687]}));
acre acre_33_38 (.clk(clk), .en(en), .top_left({trees[1637], lumberyards[1637]}), .top({trees[1638], lumberyards[1638]}), .top_right({trees[1639], lumberyards[1639]}), .left({trees[1687], lumberyards[1687]}), .right({trees[1689], lumberyards[1689]}), .bottom_left({trees[1737], lumberyards[1737]}), .bottom({trees[1738], lumberyards[1738]}), .bottom_right({trees[1739], lumberyards[1739]}), .init(2'b10), .state({trees[1688], lumberyards[1688]}));
acre acre_33_39 (.clk(clk), .en(en), .top_left({trees[1638], lumberyards[1638]}), .top({trees[1639], lumberyards[1639]}), .top_right({trees[1640], lumberyards[1640]}), .left({trees[1688], lumberyards[1688]}), .right({trees[1690], lumberyards[1690]}), .bottom_left({trees[1738], lumberyards[1738]}), .bottom({trees[1739], lumberyards[1739]}), .bottom_right({trees[1740], lumberyards[1740]}), .init(2'b01), .state({trees[1689], lumberyards[1689]}));
acre acre_33_40 (.clk(clk), .en(en), .top_left({trees[1639], lumberyards[1639]}), .top({trees[1640], lumberyards[1640]}), .top_right({trees[1641], lumberyards[1641]}), .left({trees[1689], lumberyards[1689]}), .right({trees[1691], lumberyards[1691]}), .bottom_left({trees[1739], lumberyards[1739]}), .bottom({trees[1740], lumberyards[1740]}), .bottom_right({trees[1741], lumberyards[1741]}), .init(2'b00), .state({trees[1690], lumberyards[1690]}));
acre acre_33_41 (.clk(clk), .en(en), .top_left({trees[1640], lumberyards[1640]}), .top({trees[1641], lumberyards[1641]}), .top_right({trees[1642], lumberyards[1642]}), .left({trees[1690], lumberyards[1690]}), .right({trees[1692], lumberyards[1692]}), .bottom_left({trees[1740], lumberyards[1740]}), .bottom({trees[1741], lumberyards[1741]}), .bottom_right({trees[1742], lumberyards[1742]}), .init(2'b01), .state({trees[1691], lumberyards[1691]}));
acre acre_33_42 (.clk(clk), .en(en), .top_left({trees[1641], lumberyards[1641]}), .top({trees[1642], lumberyards[1642]}), .top_right({trees[1643], lumberyards[1643]}), .left({trees[1691], lumberyards[1691]}), .right({trees[1693], lumberyards[1693]}), .bottom_left({trees[1741], lumberyards[1741]}), .bottom({trees[1742], lumberyards[1742]}), .bottom_right({trees[1743], lumberyards[1743]}), .init(2'b00), .state({trees[1692], lumberyards[1692]}));
acre acre_33_43 (.clk(clk), .en(en), .top_left({trees[1642], lumberyards[1642]}), .top({trees[1643], lumberyards[1643]}), .top_right({trees[1644], lumberyards[1644]}), .left({trees[1692], lumberyards[1692]}), .right({trees[1694], lumberyards[1694]}), .bottom_left({trees[1742], lumberyards[1742]}), .bottom({trees[1743], lumberyards[1743]}), .bottom_right({trees[1744], lumberyards[1744]}), .init(2'b00), .state({trees[1693], lumberyards[1693]}));
acre acre_33_44 (.clk(clk), .en(en), .top_left({trees[1643], lumberyards[1643]}), .top({trees[1644], lumberyards[1644]}), .top_right({trees[1645], lumberyards[1645]}), .left({trees[1693], lumberyards[1693]}), .right({trees[1695], lumberyards[1695]}), .bottom_left({trees[1743], lumberyards[1743]}), .bottom({trees[1744], lumberyards[1744]}), .bottom_right({trees[1745], lumberyards[1745]}), .init(2'b01), .state({trees[1694], lumberyards[1694]}));
acre acre_33_45 (.clk(clk), .en(en), .top_left({trees[1644], lumberyards[1644]}), .top({trees[1645], lumberyards[1645]}), .top_right({trees[1646], lumberyards[1646]}), .left({trees[1694], lumberyards[1694]}), .right({trees[1696], lumberyards[1696]}), .bottom_left({trees[1744], lumberyards[1744]}), .bottom({trees[1745], lumberyards[1745]}), .bottom_right({trees[1746], lumberyards[1746]}), .init(2'b00), .state({trees[1695], lumberyards[1695]}));
acre acre_33_46 (.clk(clk), .en(en), .top_left({trees[1645], lumberyards[1645]}), .top({trees[1646], lumberyards[1646]}), .top_right({trees[1647], lumberyards[1647]}), .left({trees[1695], lumberyards[1695]}), .right({trees[1697], lumberyards[1697]}), .bottom_left({trees[1745], lumberyards[1745]}), .bottom({trees[1746], lumberyards[1746]}), .bottom_right({trees[1747], lumberyards[1747]}), .init(2'b00), .state({trees[1696], lumberyards[1696]}));
acre acre_33_47 (.clk(clk), .en(en), .top_left({trees[1646], lumberyards[1646]}), .top({trees[1647], lumberyards[1647]}), .top_right({trees[1648], lumberyards[1648]}), .left({trees[1696], lumberyards[1696]}), .right({trees[1698], lumberyards[1698]}), .bottom_left({trees[1746], lumberyards[1746]}), .bottom({trees[1747], lumberyards[1747]}), .bottom_right({trees[1748], lumberyards[1748]}), .init(2'b10), .state({trees[1697], lumberyards[1697]}));
acre acre_33_48 (.clk(clk), .en(en), .top_left({trees[1647], lumberyards[1647]}), .top({trees[1648], lumberyards[1648]}), .top_right({trees[1649], lumberyards[1649]}), .left({trees[1697], lumberyards[1697]}), .right({trees[1699], lumberyards[1699]}), .bottom_left({trees[1747], lumberyards[1747]}), .bottom({trees[1748], lumberyards[1748]}), .bottom_right({trees[1749], lumberyards[1749]}), .init(2'b00), .state({trees[1698], lumberyards[1698]}));
acre acre_33_49 (.clk(clk), .en(en), .top_left({trees[1648], lumberyards[1648]}), .top({trees[1649], lumberyards[1649]}), .top_right(2'b0), .left({trees[1698], lumberyards[1698]}), .right(2'b0), .bottom_left({trees[1748], lumberyards[1748]}), .bottom({trees[1749], lumberyards[1749]}), .bottom_right(2'b0), .init(2'b01), .state({trees[1699], lumberyards[1699]}));
acre acre_34_0 (.clk(clk), .en(en), .top_left(2'b0), .top({trees[1650], lumberyards[1650]}), .top_right({trees[1651], lumberyards[1651]}), .left(2'b0), .right({trees[1701], lumberyards[1701]}), .bottom_left(2'b0), .bottom({trees[1750], lumberyards[1750]}), .bottom_right({trees[1751], lumberyards[1751]}), .init(2'b10), .state({trees[1700], lumberyards[1700]}));
acre acre_34_1 (.clk(clk), .en(en), .top_left({trees[1650], lumberyards[1650]}), .top({trees[1651], lumberyards[1651]}), .top_right({trees[1652], lumberyards[1652]}), .left({trees[1700], lumberyards[1700]}), .right({trees[1702], lumberyards[1702]}), .bottom_left({trees[1750], lumberyards[1750]}), .bottom({trees[1751], lumberyards[1751]}), .bottom_right({trees[1752], lumberyards[1752]}), .init(2'b00), .state({trees[1701], lumberyards[1701]}));
acre acre_34_2 (.clk(clk), .en(en), .top_left({trees[1651], lumberyards[1651]}), .top({trees[1652], lumberyards[1652]}), .top_right({trees[1653], lumberyards[1653]}), .left({trees[1701], lumberyards[1701]}), .right({trees[1703], lumberyards[1703]}), .bottom_left({trees[1751], lumberyards[1751]}), .bottom({trees[1752], lumberyards[1752]}), .bottom_right({trees[1753], lumberyards[1753]}), .init(2'b10), .state({trees[1702], lumberyards[1702]}));
acre acre_34_3 (.clk(clk), .en(en), .top_left({trees[1652], lumberyards[1652]}), .top({trees[1653], lumberyards[1653]}), .top_right({trees[1654], lumberyards[1654]}), .left({trees[1702], lumberyards[1702]}), .right({trees[1704], lumberyards[1704]}), .bottom_left({trees[1752], lumberyards[1752]}), .bottom({trees[1753], lumberyards[1753]}), .bottom_right({trees[1754], lumberyards[1754]}), .init(2'b00), .state({trees[1703], lumberyards[1703]}));
acre acre_34_4 (.clk(clk), .en(en), .top_left({trees[1653], lumberyards[1653]}), .top({trees[1654], lumberyards[1654]}), .top_right({trees[1655], lumberyards[1655]}), .left({trees[1703], lumberyards[1703]}), .right({trees[1705], lumberyards[1705]}), .bottom_left({trees[1753], lumberyards[1753]}), .bottom({trees[1754], lumberyards[1754]}), .bottom_right({trees[1755], lumberyards[1755]}), .init(2'b00), .state({trees[1704], lumberyards[1704]}));
acre acre_34_5 (.clk(clk), .en(en), .top_left({trees[1654], lumberyards[1654]}), .top({trees[1655], lumberyards[1655]}), .top_right({trees[1656], lumberyards[1656]}), .left({trees[1704], lumberyards[1704]}), .right({trees[1706], lumberyards[1706]}), .bottom_left({trees[1754], lumberyards[1754]}), .bottom({trees[1755], lumberyards[1755]}), .bottom_right({trees[1756], lumberyards[1756]}), .init(2'b00), .state({trees[1705], lumberyards[1705]}));
acre acre_34_6 (.clk(clk), .en(en), .top_left({trees[1655], lumberyards[1655]}), .top({trees[1656], lumberyards[1656]}), .top_right({trees[1657], lumberyards[1657]}), .left({trees[1705], lumberyards[1705]}), .right({trees[1707], lumberyards[1707]}), .bottom_left({trees[1755], lumberyards[1755]}), .bottom({trees[1756], lumberyards[1756]}), .bottom_right({trees[1757], lumberyards[1757]}), .init(2'b00), .state({trees[1706], lumberyards[1706]}));
acre acre_34_7 (.clk(clk), .en(en), .top_left({trees[1656], lumberyards[1656]}), .top({trees[1657], lumberyards[1657]}), .top_right({trees[1658], lumberyards[1658]}), .left({trees[1706], lumberyards[1706]}), .right({trees[1708], lumberyards[1708]}), .bottom_left({trees[1756], lumberyards[1756]}), .bottom({trees[1757], lumberyards[1757]}), .bottom_right({trees[1758], lumberyards[1758]}), .init(2'b00), .state({trees[1707], lumberyards[1707]}));
acre acre_34_8 (.clk(clk), .en(en), .top_left({trees[1657], lumberyards[1657]}), .top({trees[1658], lumberyards[1658]}), .top_right({trees[1659], lumberyards[1659]}), .left({trees[1707], lumberyards[1707]}), .right({trees[1709], lumberyards[1709]}), .bottom_left({trees[1757], lumberyards[1757]}), .bottom({trees[1758], lumberyards[1758]}), .bottom_right({trees[1759], lumberyards[1759]}), .init(2'b00), .state({trees[1708], lumberyards[1708]}));
acre acre_34_9 (.clk(clk), .en(en), .top_left({trees[1658], lumberyards[1658]}), .top({trees[1659], lumberyards[1659]}), .top_right({trees[1660], lumberyards[1660]}), .left({trees[1708], lumberyards[1708]}), .right({trees[1710], lumberyards[1710]}), .bottom_left({trees[1758], lumberyards[1758]}), .bottom({trees[1759], lumberyards[1759]}), .bottom_right({trees[1760], lumberyards[1760]}), .init(2'b10), .state({trees[1709], lumberyards[1709]}));
acre acre_34_10 (.clk(clk), .en(en), .top_left({trees[1659], lumberyards[1659]}), .top({trees[1660], lumberyards[1660]}), .top_right({trees[1661], lumberyards[1661]}), .left({trees[1709], lumberyards[1709]}), .right({trees[1711], lumberyards[1711]}), .bottom_left({trees[1759], lumberyards[1759]}), .bottom({trees[1760], lumberyards[1760]}), .bottom_right({trees[1761], lumberyards[1761]}), .init(2'b00), .state({trees[1710], lumberyards[1710]}));
acre acre_34_11 (.clk(clk), .en(en), .top_left({trees[1660], lumberyards[1660]}), .top({trees[1661], lumberyards[1661]}), .top_right({trees[1662], lumberyards[1662]}), .left({trees[1710], lumberyards[1710]}), .right({trees[1712], lumberyards[1712]}), .bottom_left({trees[1760], lumberyards[1760]}), .bottom({trees[1761], lumberyards[1761]}), .bottom_right({trees[1762], lumberyards[1762]}), .init(2'b10), .state({trees[1711], lumberyards[1711]}));
acre acre_34_12 (.clk(clk), .en(en), .top_left({trees[1661], lumberyards[1661]}), .top({trees[1662], lumberyards[1662]}), .top_right({trees[1663], lumberyards[1663]}), .left({trees[1711], lumberyards[1711]}), .right({trees[1713], lumberyards[1713]}), .bottom_left({trees[1761], lumberyards[1761]}), .bottom({trees[1762], lumberyards[1762]}), .bottom_right({trees[1763], lumberyards[1763]}), .init(2'b01), .state({trees[1712], lumberyards[1712]}));
acre acre_34_13 (.clk(clk), .en(en), .top_left({trees[1662], lumberyards[1662]}), .top({trees[1663], lumberyards[1663]}), .top_right({trees[1664], lumberyards[1664]}), .left({trees[1712], lumberyards[1712]}), .right({trees[1714], lumberyards[1714]}), .bottom_left({trees[1762], lumberyards[1762]}), .bottom({trees[1763], lumberyards[1763]}), .bottom_right({trees[1764], lumberyards[1764]}), .init(2'b00), .state({trees[1713], lumberyards[1713]}));
acre acre_34_14 (.clk(clk), .en(en), .top_left({trees[1663], lumberyards[1663]}), .top({trees[1664], lumberyards[1664]}), .top_right({trees[1665], lumberyards[1665]}), .left({trees[1713], lumberyards[1713]}), .right({trees[1715], lumberyards[1715]}), .bottom_left({trees[1763], lumberyards[1763]}), .bottom({trees[1764], lumberyards[1764]}), .bottom_right({trees[1765], lumberyards[1765]}), .init(2'b00), .state({trees[1714], lumberyards[1714]}));
acre acre_34_15 (.clk(clk), .en(en), .top_left({trees[1664], lumberyards[1664]}), .top({trees[1665], lumberyards[1665]}), .top_right({trees[1666], lumberyards[1666]}), .left({trees[1714], lumberyards[1714]}), .right({trees[1716], lumberyards[1716]}), .bottom_left({trees[1764], lumberyards[1764]}), .bottom({trees[1765], lumberyards[1765]}), .bottom_right({trees[1766], lumberyards[1766]}), .init(2'b00), .state({trees[1715], lumberyards[1715]}));
acre acre_34_16 (.clk(clk), .en(en), .top_left({trees[1665], lumberyards[1665]}), .top({trees[1666], lumberyards[1666]}), .top_right({trees[1667], lumberyards[1667]}), .left({trees[1715], lumberyards[1715]}), .right({trees[1717], lumberyards[1717]}), .bottom_left({trees[1765], lumberyards[1765]}), .bottom({trees[1766], lumberyards[1766]}), .bottom_right({trees[1767], lumberyards[1767]}), .init(2'b00), .state({trees[1716], lumberyards[1716]}));
acre acre_34_17 (.clk(clk), .en(en), .top_left({trees[1666], lumberyards[1666]}), .top({trees[1667], lumberyards[1667]}), .top_right({trees[1668], lumberyards[1668]}), .left({trees[1716], lumberyards[1716]}), .right({trees[1718], lumberyards[1718]}), .bottom_left({trees[1766], lumberyards[1766]}), .bottom({trees[1767], lumberyards[1767]}), .bottom_right({trees[1768], lumberyards[1768]}), .init(2'b01), .state({trees[1717], lumberyards[1717]}));
acre acre_34_18 (.clk(clk), .en(en), .top_left({trees[1667], lumberyards[1667]}), .top({trees[1668], lumberyards[1668]}), .top_right({trees[1669], lumberyards[1669]}), .left({trees[1717], lumberyards[1717]}), .right({trees[1719], lumberyards[1719]}), .bottom_left({trees[1767], lumberyards[1767]}), .bottom({trees[1768], lumberyards[1768]}), .bottom_right({trees[1769], lumberyards[1769]}), .init(2'b01), .state({trees[1718], lumberyards[1718]}));
acre acre_34_19 (.clk(clk), .en(en), .top_left({trees[1668], lumberyards[1668]}), .top({trees[1669], lumberyards[1669]}), .top_right({trees[1670], lumberyards[1670]}), .left({trees[1718], lumberyards[1718]}), .right({trees[1720], lumberyards[1720]}), .bottom_left({trees[1768], lumberyards[1768]}), .bottom({trees[1769], lumberyards[1769]}), .bottom_right({trees[1770], lumberyards[1770]}), .init(2'b10), .state({trees[1719], lumberyards[1719]}));
acre acre_34_20 (.clk(clk), .en(en), .top_left({trees[1669], lumberyards[1669]}), .top({trees[1670], lumberyards[1670]}), .top_right({trees[1671], lumberyards[1671]}), .left({trees[1719], lumberyards[1719]}), .right({trees[1721], lumberyards[1721]}), .bottom_left({trees[1769], lumberyards[1769]}), .bottom({trees[1770], lumberyards[1770]}), .bottom_right({trees[1771], lumberyards[1771]}), .init(2'b10), .state({trees[1720], lumberyards[1720]}));
acre acre_34_21 (.clk(clk), .en(en), .top_left({trees[1670], lumberyards[1670]}), .top({trees[1671], lumberyards[1671]}), .top_right({trees[1672], lumberyards[1672]}), .left({trees[1720], lumberyards[1720]}), .right({trees[1722], lumberyards[1722]}), .bottom_left({trees[1770], lumberyards[1770]}), .bottom({trees[1771], lumberyards[1771]}), .bottom_right({trees[1772], lumberyards[1772]}), .init(2'b01), .state({trees[1721], lumberyards[1721]}));
acre acre_34_22 (.clk(clk), .en(en), .top_left({trees[1671], lumberyards[1671]}), .top({trees[1672], lumberyards[1672]}), .top_right({trees[1673], lumberyards[1673]}), .left({trees[1721], lumberyards[1721]}), .right({trees[1723], lumberyards[1723]}), .bottom_left({trees[1771], lumberyards[1771]}), .bottom({trees[1772], lumberyards[1772]}), .bottom_right({trees[1773], lumberyards[1773]}), .init(2'b00), .state({trees[1722], lumberyards[1722]}));
acre acre_34_23 (.clk(clk), .en(en), .top_left({trees[1672], lumberyards[1672]}), .top({trees[1673], lumberyards[1673]}), .top_right({trees[1674], lumberyards[1674]}), .left({trees[1722], lumberyards[1722]}), .right({trees[1724], lumberyards[1724]}), .bottom_left({trees[1772], lumberyards[1772]}), .bottom({trees[1773], lumberyards[1773]}), .bottom_right({trees[1774], lumberyards[1774]}), .init(2'b00), .state({trees[1723], lumberyards[1723]}));
acre acre_34_24 (.clk(clk), .en(en), .top_left({trees[1673], lumberyards[1673]}), .top({trees[1674], lumberyards[1674]}), .top_right({trees[1675], lumberyards[1675]}), .left({trees[1723], lumberyards[1723]}), .right({trees[1725], lumberyards[1725]}), .bottom_left({trees[1773], lumberyards[1773]}), .bottom({trees[1774], lumberyards[1774]}), .bottom_right({trees[1775], lumberyards[1775]}), .init(2'b10), .state({trees[1724], lumberyards[1724]}));
acre acre_34_25 (.clk(clk), .en(en), .top_left({trees[1674], lumberyards[1674]}), .top({trees[1675], lumberyards[1675]}), .top_right({trees[1676], lumberyards[1676]}), .left({trees[1724], lumberyards[1724]}), .right({trees[1726], lumberyards[1726]}), .bottom_left({trees[1774], lumberyards[1774]}), .bottom({trees[1775], lumberyards[1775]}), .bottom_right({trees[1776], lumberyards[1776]}), .init(2'b00), .state({trees[1725], lumberyards[1725]}));
acre acre_34_26 (.clk(clk), .en(en), .top_left({trees[1675], lumberyards[1675]}), .top({trees[1676], lumberyards[1676]}), .top_right({trees[1677], lumberyards[1677]}), .left({trees[1725], lumberyards[1725]}), .right({trees[1727], lumberyards[1727]}), .bottom_left({trees[1775], lumberyards[1775]}), .bottom({trees[1776], lumberyards[1776]}), .bottom_right({trees[1777], lumberyards[1777]}), .init(2'b00), .state({trees[1726], lumberyards[1726]}));
acre acre_34_27 (.clk(clk), .en(en), .top_left({trees[1676], lumberyards[1676]}), .top({trees[1677], lumberyards[1677]}), .top_right({trees[1678], lumberyards[1678]}), .left({trees[1726], lumberyards[1726]}), .right({trees[1728], lumberyards[1728]}), .bottom_left({trees[1776], lumberyards[1776]}), .bottom({trees[1777], lumberyards[1777]}), .bottom_right({trees[1778], lumberyards[1778]}), .init(2'b01), .state({trees[1727], lumberyards[1727]}));
acre acre_34_28 (.clk(clk), .en(en), .top_left({trees[1677], lumberyards[1677]}), .top({trees[1678], lumberyards[1678]}), .top_right({trees[1679], lumberyards[1679]}), .left({trees[1727], lumberyards[1727]}), .right({trees[1729], lumberyards[1729]}), .bottom_left({trees[1777], lumberyards[1777]}), .bottom({trees[1778], lumberyards[1778]}), .bottom_right({trees[1779], lumberyards[1779]}), .init(2'b10), .state({trees[1728], lumberyards[1728]}));
acre acre_34_29 (.clk(clk), .en(en), .top_left({trees[1678], lumberyards[1678]}), .top({trees[1679], lumberyards[1679]}), .top_right({trees[1680], lumberyards[1680]}), .left({trees[1728], lumberyards[1728]}), .right({trees[1730], lumberyards[1730]}), .bottom_left({trees[1778], lumberyards[1778]}), .bottom({trees[1779], lumberyards[1779]}), .bottom_right({trees[1780], lumberyards[1780]}), .init(2'b00), .state({trees[1729], lumberyards[1729]}));
acre acre_34_30 (.clk(clk), .en(en), .top_left({trees[1679], lumberyards[1679]}), .top({trees[1680], lumberyards[1680]}), .top_right({trees[1681], lumberyards[1681]}), .left({trees[1729], lumberyards[1729]}), .right({trees[1731], lumberyards[1731]}), .bottom_left({trees[1779], lumberyards[1779]}), .bottom({trees[1780], lumberyards[1780]}), .bottom_right({trees[1781], lumberyards[1781]}), .init(2'b00), .state({trees[1730], lumberyards[1730]}));
acre acre_34_31 (.clk(clk), .en(en), .top_left({trees[1680], lumberyards[1680]}), .top({trees[1681], lumberyards[1681]}), .top_right({trees[1682], lumberyards[1682]}), .left({trees[1730], lumberyards[1730]}), .right({trees[1732], lumberyards[1732]}), .bottom_left({trees[1780], lumberyards[1780]}), .bottom({trees[1781], lumberyards[1781]}), .bottom_right({trees[1782], lumberyards[1782]}), .init(2'b00), .state({trees[1731], lumberyards[1731]}));
acre acre_34_32 (.clk(clk), .en(en), .top_left({trees[1681], lumberyards[1681]}), .top({trees[1682], lumberyards[1682]}), .top_right({trees[1683], lumberyards[1683]}), .left({trees[1731], lumberyards[1731]}), .right({trees[1733], lumberyards[1733]}), .bottom_left({trees[1781], lumberyards[1781]}), .bottom({trees[1782], lumberyards[1782]}), .bottom_right({trees[1783], lumberyards[1783]}), .init(2'b00), .state({trees[1732], lumberyards[1732]}));
acre acre_34_33 (.clk(clk), .en(en), .top_left({trees[1682], lumberyards[1682]}), .top({trees[1683], lumberyards[1683]}), .top_right({trees[1684], lumberyards[1684]}), .left({trees[1732], lumberyards[1732]}), .right({trees[1734], lumberyards[1734]}), .bottom_left({trees[1782], lumberyards[1782]}), .bottom({trees[1783], lumberyards[1783]}), .bottom_right({trees[1784], lumberyards[1784]}), .init(2'b10), .state({trees[1733], lumberyards[1733]}));
acre acre_34_34 (.clk(clk), .en(en), .top_left({trees[1683], lumberyards[1683]}), .top({trees[1684], lumberyards[1684]}), .top_right({trees[1685], lumberyards[1685]}), .left({trees[1733], lumberyards[1733]}), .right({trees[1735], lumberyards[1735]}), .bottom_left({trees[1783], lumberyards[1783]}), .bottom({trees[1784], lumberyards[1784]}), .bottom_right({trees[1785], lumberyards[1785]}), .init(2'b10), .state({trees[1734], lumberyards[1734]}));
acre acre_34_35 (.clk(clk), .en(en), .top_left({trees[1684], lumberyards[1684]}), .top({trees[1685], lumberyards[1685]}), .top_right({trees[1686], lumberyards[1686]}), .left({trees[1734], lumberyards[1734]}), .right({trees[1736], lumberyards[1736]}), .bottom_left({trees[1784], lumberyards[1784]}), .bottom({trees[1785], lumberyards[1785]}), .bottom_right({trees[1786], lumberyards[1786]}), .init(2'b10), .state({trees[1735], lumberyards[1735]}));
acre acre_34_36 (.clk(clk), .en(en), .top_left({trees[1685], lumberyards[1685]}), .top({trees[1686], lumberyards[1686]}), .top_right({trees[1687], lumberyards[1687]}), .left({trees[1735], lumberyards[1735]}), .right({trees[1737], lumberyards[1737]}), .bottom_left({trees[1785], lumberyards[1785]}), .bottom({trees[1786], lumberyards[1786]}), .bottom_right({trees[1787], lumberyards[1787]}), .init(2'b10), .state({trees[1736], lumberyards[1736]}));
acre acre_34_37 (.clk(clk), .en(en), .top_left({trees[1686], lumberyards[1686]}), .top({trees[1687], lumberyards[1687]}), .top_right({trees[1688], lumberyards[1688]}), .left({trees[1736], lumberyards[1736]}), .right({trees[1738], lumberyards[1738]}), .bottom_left({trees[1786], lumberyards[1786]}), .bottom({trees[1787], lumberyards[1787]}), .bottom_right({trees[1788], lumberyards[1788]}), .init(2'b00), .state({trees[1737], lumberyards[1737]}));
acre acre_34_38 (.clk(clk), .en(en), .top_left({trees[1687], lumberyards[1687]}), .top({trees[1688], lumberyards[1688]}), .top_right({trees[1689], lumberyards[1689]}), .left({trees[1737], lumberyards[1737]}), .right({trees[1739], lumberyards[1739]}), .bottom_left({trees[1787], lumberyards[1787]}), .bottom({trees[1788], lumberyards[1788]}), .bottom_right({trees[1789], lumberyards[1789]}), .init(2'b10), .state({trees[1738], lumberyards[1738]}));
acre acre_34_39 (.clk(clk), .en(en), .top_left({trees[1688], lumberyards[1688]}), .top({trees[1689], lumberyards[1689]}), .top_right({trees[1690], lumberyards[1690]}), .left({trees[1738], lumberyards[1738]}), .right({trees[1740], lumberyards[1740]}), .bottom_left({trees[1788], lumberyards[1788]}), .bottom({trees[1789], lumberyards[1789]}), .bottom_right({trees[1790], lumberyards[1790]}), .init(2'b10), .state({trees[1739], lumberyards[1739]}));
acre acre_34_40 (.clk(clk), .en(en), .top_left({trees[1689], lumberyards[1689]}), .top({trees[1690], lumberyards[1690]}), .top_right({trees[1691], lumberyards[1691]}), .left({trees[1739], lumberyards[1739]}), .right({trees[1741], lumberyards[1741]}), .bottom_left({trees[1789], lumberyards[1789]}), .bottom({trees[1790], lumberyards[1790]}), .bottom_right({trees[1791], lumberyards[1791]}), .init(2'b00), .state({trees[1740], lumberyards[1740]}));
acre acre_34_41 (.clk(clk), .en(en), .top_left({trees[1690], lumberyards[1690]}), .top({trees[1691], lumberyards[1691]}), .top_right({trees[1692], lumberyards[1692]}), .left({trees[1740], lumberyards[1740]}), .right({trees[1742], lumberyards[1742]}), .bottom_left({trees[1790], lumberyards[1790]}), .bottom({trees[1791], lumberyards[1791]}), .bottom_right({trees[1792], lumberyards[1792]}), .init(2'b00), .state({trees[1741], lumberyards[1741]}));
acre acre_34_42 (.clk(clk), .en(en), .top_left({trees[1691], lumberyards[1691]}), .top({trees[1692], lumberyards[1692]}), .top_right({trees[1693], lumberyards[1693]}), .left({trees[1741], lumberyards[1741]}), .right({trees[1743], lumberyards[1743]}), .bottom_left({trees[1791], lumberyards[1791]}), .bottom({trees[1792], lumberyards[1792]}), .bottom_right({trees[1793], lumberyards[1793]}), .init(2'b01), .state({trees[1742], lumberyards[1742]}));
acre acre_34_43 (.clk(clk), .en(en), .top_left({trees[1692], lumberyards[1692]}), .top({trees[1693], lumberyards[1693]}), .top_right({trees[1694], lumberyards[1694]}), .left({trees[1742], lumberyards[1742]}), .right({trees[1744], lumberyards[1744]}), .bottom_left({trees[1792], lumberyards[1792]}), .bottom({trees[1793], lumberyards[1793]}), .bottom_right({trees[1794], lumberyards[1794]}), .init(2'b00), .state({trees[1743], lumberyards[1743]}));
acre acre_34_44 (.clk(clk), .en(en), .top_left({trees[1693], lumberyards[1693]}), .top({trees[1694], lumberyards[1694]}), .top_right({trees[1695], lumberyards[1695]}), .left({trees[1743], lumberyards[1743]}), .right({trees[1745], lumberyards[1745]}), .bottom_left({trees[1793], lumberyards[1793]}), .bottom({trees[1794], lumberyards[1794]}), .bottom_right({trees[1795], lumberyards[1795]}), .init(2'b00), .state({trees[1744], lumberyards[1744]}));
acre acre_34_45 (.clk(clk), .en(en), .top_left({trees[1694], lumberyards[1694]}), .top({trees[1695], lumberyards[1695]}), .top_right({trees[1696], lumberyards[1696]}), .left({trees[1744], lumberyards[1744]}), .right({trees[1746], lumberyards[1746]}), .bottom_left({trees[1794], lumberyards[1794]}), .bottom({trees[1795], lumberyards[1795]}), .bottom_right({trees[1796], lumberyards[1796]}), .init(2'b00), .state({trees[1745], lumberyards[1745]}));
acre acre_34_46 (.clk(clk), .en(en), .top_left({trees[1695], lumberyards[1695]}), .top({trees[1696], lumberyards[1696]}), .top_right({trees[1697], lumberyards[1697]}), .left({trees[1745], lumberyards[1745]}), .right({trees[1747], lumberyards[1747]}), .bottom_left({trees[1795], lumberyards[1795]}), .bottom({trees[1796], lumberyards[1796]}), .bottom_right({trees[1797], lumberyards[1797]}), .init(2'b00), .state({trees[1746], lumberyards[1746]}));
acre acre_34_47 (.clk(clk), .en(en), .top_left({trees[1696], lumberyards[1696]}), .top({trees[1697], lumberyards[1697]}), .top_right({trees[1698], lumberyards[1698]}), .left({trees[1746], lumberyards[1746]}), .right({trees[1748], lumberyards[1748]}), .bottom_left({trees[1796], lumberyards[1796]}), .bottom({trees[1797], lumberyards[1797]}), .bottom_right({trees[1798], lumberyards[1798]}), .init(2'b01), .state({trees[1747], lumberyards[1747]}));
acre acre_34_48 (.clk(clk), .en(en), .top_left({trees[1697], lumberyards[1697]}), .top({trees[1698], lumberyards[1698]}), .top_right({trees[1699], lumberyards[1699]}), .left({trees[1747], lumberyards[1747]}), .right({trees[1749], lumberyards[1749]}), .bottom_left({trees[1797], lumberyards[1797]}), .bottom({trees[1798], lumberyards[1798]}), .bottom_right({trees[1799], lumberyards[1799]}), .init(2'b00), .state({trees[1748], lumberyards[1748]}));
acre acre_34_49 (.clk(clk), .en(en), .top_left({trees[1698], lumberyards[1698]}), .top({trees[1699], lumberyards[1699]}), .top_right(2'b0), .left({trees[1748], lumberyards[1748]}), .right(2'b0), .bottom_left({trees[1798], lumberyards[1798]}), .bottom({trees[1799], lumberyards[1799]}), .bottom_right(2'b0), .init(2'b10), .state({trees[1749], lumberyards[1749]}));
acre acre_35_0 (.clk(clk), .en(en), .top_left(2'b0), .top({trees[1700], lumberyards[1700]}), .top_right({trees[1701], lumberyards[1701]}), .left(2'b0), .right({trees[1751], lumberyards[1751]}), .bottom_left(2'b0), .bottom({trees[1800], lumberyards[1800]}), .bottom_right({trees[1801], lumberyards[1801]}), .init(2'b00), .state({trees[1750], lumberyards[1750]}));
acre acre_35_1 (.clk(clk), .en(en), .top_left({trees[1700], lumberyards[1700]}), .top({trees[1701], lumberyards[1701]}), .top_right({trees[1702], lumberyards[1702]}), .left({trees[1750], lumberyards[1750]}), .right({trees[1752], lumberyards[1752]}), .bottom_left({trees[1800], lumberyards[1800]}), .bottom({trees[1801], lumberyards[1801]}), .bottom_right({trees[1802], lumberyards[1802]}), .init(2'b10), .state({trees[1751], lumberyards[1751]}));
acre acre_35_2 (.clk(clk), .en(en), .top_left({trees[1701], lumberyards[1701]}), .top({trees[1702], lumberyards[1702]}), .top_right({trees[1703], lumberyards[1703]}), .left({trees[1751], lumberyards[1751]}), .right({trees[1753], lumberyards[1753]}), .bottom_left({trees[1801], lumberyards[1801]}), .bottom({trees[1802], lumberyards[1802]}), .bottom_right({trees[1803], lumberyards[1803]}), .init(2'b00), .state({trees[1752], lumberyards[1752]}));
acre acre_35_3 (.clk(clk), .en(en), .top_left({trees[1702], lumberyards[1702]}), .top({trees[1703], lumberyards[1703]}), .top_right({trees[1704], lumberyards[1704]}), .left({trees[1752], lumberyards[1752]}), .right({trees[1754], lumberyards[1754]}), .bottom_left({trees[1802], lumberyards[1802]}), .bottom({trees[1803], lumberyards[1803]}), .bottom_right({trees[1804], lumberyards[1804]}), .init(2'b00), .state({trees[1753], lumberyards[1753]}));
acre acre_35_4 (.clk(clk), .en(en), .top_left({trees[1703], lumberyards[1703]}), .top({trees[1704], lumberyards[1704]}), .top_right({trees[1705], lumberyards[1705]}), .left({trees[1753], lumberyards[1753]}), .right({trees[1755], lumberyards[1755]}), .bottom_left({trees[1803], lumberyards[1803]}), .bottom({trees[1804], lumberyards[1804]}), .bottom_right({trees[1805], lumberyards[1805]}), .init(2'b01), .state({trees[1754], lumberyards[1754]}));
acre acre_35_5 (.clk(clk), .en(en), .top_left({trees[1704], lumberyards[1704]}), .top({trees[1705], lumberyards[1705]}), .top_right({trees[1706], lumberyards[1706]}), .left({trees[1754], lumberyards[1754]}), .right({trees[1756], lumberyards[1756]}), .bottom_left({trees[1804], lumberyards[1804]}), .bottom({trees[1805], lumberyards[1805]}), .bottom_right({trees[1806], lumberyards[1806]}), .init(2'b10), .state({trees[1755], lumberyards[1755]}));
acre acre_35_6 (.clk(clk), .en(en), .top_left({trees[1705], lumberyards[1705]}), .top({trees[1706], lumberyards[1706]}), .top_right({trees[1707], lumberyards[1707]}), .left({trees[1755], lumberyards[1755]}), .right({trees[1757], lumberyards[1757]}), .bottom_left({trees[1805], lumberyards[1805]}), .bottom({trees[1806], lumberyards[1806]}), .bottom_right({trees[1807], lumberyards[1807]}), .init(2'b01), .state({trees[1756], lumberyards[1756]}));
acre acre_35_7 (.clk(clk), .en(en), .top_left({trees[1706], lumberyards[1706]}), .top({trees[1707], lumberyards[1707]}), .top_right({trees[1708], lumberyards[1708]}), .left({trees[1756], lumberyards[1756]}), .right({trees[1758], lumberyards[1758]}), .bottom_left({trees[1806], lumberyards[1806]}), .bottom({trees[1807], lumberyards[1807]}), .bottom_right({trees[1808], lumberyards[1808]}), .init(2'b00), .state({trees[1757], lumberyards[1757]}));
acre acre_35_8 (.clk(clk), .en(en), .top_left({trees[1707], lumberyards[1707]}), .top({trees[1708], lumberyards[1708]}), .top_right({trees[1709], lumberyards[1709]}), .left({trees[1757], lumberyards[1757]}), .right({trees[1759], lumberyards[1759]}), .bottom_left({trees[1807], lumberyards[1807]}), .bottom({trees[1808], lumberyards[1808]}), .bottom_right({trees[1809], lumberyards[1809]}), .init(2'b00), .state({trees[1758], lumberyards[1758]}));
acre acre_35_9 (.clk(clk), .en(en), .top_left({trees[1708], lumberyards[1708]}), .top({trees[1709], lumberyards[1709]}), .top_right({trees[1710], lumberyards[1710]}), .left({trees[1758], lumberyards[1758]}), .right({trees[1760], lumberyards[1760]}), .bottom_left({trees[1808], lumberyards[1808]}), .bottom({trees[1809], lumberyards[1809]}), .bottom_right({trees[1810], lumberyards[1810]}), .init(2'b10), .state({trees[1759], lumberyards[1759]}));
acre acre_35_10 (.clk(clk), .en(en), .top_left({trees[1709], lumberyards[1709]}), .top({trees[1710], lumberyards[1710]}), .top_right({trees[1711], lumberyards[1711]}), .left({trees[1759], lumberyards[1759]}), .right({trees[1761], lumberyards[1761]}), .bottom_left({trees[1809], lumberyards[1809]}), .bottom({trees[1810], lumberyards[1810]}), .bottom_right({trees[1811], lumberyards[1811]}), .init(2'b00), .state({trees[1760], lumberyards[1760]}));
acre acre_35_11 (.clk(clk), .en(en), .top_left({trees[1710], lumberyards[1710]}), .top({trees[1711], lumberyards[1711]}), .top_right({trees[1712], lumberyards[1712]}), .left({trees[1760], lumberyards[1760]}), .right({trees[1762], lumberyards[1762]}), .bottom_left({trees[1810], lumberyards[1810]}), .bottom({trees[1811], lumberyards[1811]}), .bottom_right({trees[1812], lumberyards[1812]}), .init(2'b00), .state({trees[1761], lumberyards[1761]}));
acre acre_35_12 (.clk(clk), .en(en), .top_left({trees[1711], lumberyards[1711]}), .top({trees[1712], lumberyards[1712]}), .top_right({trees[1713], lumberyards[1713]}), .left({trees[1761], lumberyards[1761]}), .right({trees[1763], lumberyards[1763]}), .bottom_left({trees[1811], lumberyards[1811]}), .bottom({trees[1812], lumberyards[1812]}), .bottom_right({trees[1813], lumberyards[1813]}), .init(2'b01), .state({trees[1762], lumberyards[1762]}));
acre acre_35_13 (.clk(clk), .en(en), .top_left({trees[1712], lumberyards[1712]}), .top({trees[1713], lumberyards[1713]}), .top_right({trees[1714], lumberyards[1714]}), .left({trees[1762], lumberyards[1762]}), .right({trees[1764], lumberyards[1764]}), .bottom_left({trees[1812], lumberyards[1812]}), .bottom({trees[1813], lumberyards[1813]}), .bottom_right({trees[1814], lumberyards[1814]}), .init(2'b01), .state({trees[1763], lumberyards[1763]}));
acre acre_35_14 (.clk(clk), .en(en), .top_left({trees[1713], lumberyards[1713]}), .top({trees[1714], lumberyards[1714]}), .top_right({trees[1715], lumberyards[1715]}), .left({trees[1763], lumberyards[1763]}), .right({trees[1765], lumberyards[1765]}), .bottom_left({trees[1813], lumberyards[1813]}), .bottom({trees[1814], lumberyards[1814]}), .bottom_right({trees[1815], lumberyards[1815]}), .init(2'b10), .state({trees[1764], lumberyards[1764]}));
acre acre_35_15 (.clk(clk), .en(en), .top_left({trees[1714], lumberyards[1714]}), .top({trees[1715], lumberyards[1715]}), .top_right({trees[1716], lumberyards[1716]}), .left({trees[1764], lumberyards[1764]}), .right({trees[1766], lumberyards[1766]}), .bottom_left({trees[1814], lumberyards[1814]}), .bottom({trees[1815], lumberyards[1815]}), .bottom_right({trees[1816], lumberyards[1816]}), .init(2'b10), .state({trees[1765], lumberyards[1765]}));
acre acre_35_16 (.clk(clk), .en(en), .top_left({trees[1715], lumberyards[1715]}), .top({trees[1716], lumberyards[1716]}), .top_right({trees[1717], lumberyards[1717]}), .left({trees[1765], lumberyards[1765]}), .right({trees[1767], lumberyards[1767]}), .bottom_left({trees[1815], lumberyards[1815]}), .bottom({trees[1816], lumberyards[1816]}), .bottom_right({trees[1817], lumberyards[1817]}), .init(2'b01), .state({trees[1766], lumberyards[1766]}));
acre acre_35_17 (.clk(clk), .en(en), .top_left({trees[1716], lumberyards[1716]}), .top({trees[1717], lumberyards[1717]}), .top_right({trees[1718], lumberyards[1718]}), .left({trees[1766], lumberyards[1766]}), .right({trees[1768], lumberyards[1768]}), .bottom_left({trees[1816], lumberyards[1816]}), .bottom({trees[1817], lumberyards[1817]}), .bottom_right({trees[1818], lumberyards[1818]}), .init(2'b00), .state({trees[1767], lumberyards[1767]}));
acre acre_35_18 (.clk(clk), .en(en), .top_left({trees[1717], lumberyards[1717]}), .top({trees[1718], lumberyards[1718]}), .top_right({trees[1719], lumberyards[1719]}), .left({trees[1767], lumberyards[1767]}), .right({trees[1769], lumberyards[1769]}), .bottom_left({trees[1817], lumberyards[1817]}), .bottom({trees[1818], lumberyards[1818]}), .bottom_right({trees[1819], lumberyards[1819]}), .init(2'b01), .state({trees[1768], lumberyards[1768]}));
acre acre_35_19 (.clk(clk), .en(en), .top_left({trees[1718], lumberyards[1718]}), .top({trees[1719], lumberyards[1719]}), .top_right({trees[1720], lumberyards[1720]}), .left({trees[1768], lumberyards[1768]}), .right({trees[1770], lumberyards[1770]}), .bottom_left({trees[1818], lumberyards[1818]}), .bottom({trees[1819], lumberyards[1819]}), .bottom_right({trees[1820], lumberyards[1820]}), .init(2'b00), .state({trees[1769], lumberyards[1769]}));
acre acre_35_20 (.clk(clk), .en(en), .top_left({trees[1719], lumberyards[1719]}), .top({trees[1720], lumberyards[1720]}), .top_right({trees[1721], lumberyards[1721]}), .left({trees[1769], lumberyards[1769]}), .right({trees[1771], lumberyards[1771]}), .bottom_left({trees[1819], lumberyards[1819]}), .bottom({trees[1820], lumberyards[1820]}), .bottom_right({trees[1821], lumberyards[1821]}), .init(2'b10), .state({trees[1770], lumberyards[1770]}));
acre acre_35_21 (.clk(clk), .en(en), .top_left({trees[1720], lumberyards[1720]}), .top({trees[1721], lumberyards[1721]}), .top_right({trees[1722], lumberyards[1722]}), .left({trees[1770], lumberyards[1770]}), .right({trees[1772], lumberyards[1772]}), .bottom_left({trees[1820], lumberyards[1820]}), .bottom({trees[1821], lumberyards[1821]}), .bottom_right({trees[1822], lumberyards[1822]}), .init(2'b00), .state({trees[1771], lumberyards[1771]}));
acre acre_35_22 (.clk(clk), .en(en), .top_left({trees[1721], lumberyards[1721]}), .top({trees[1722], lumberyards[1722]}), .top_right({trees[1723], lumberyards[1723]}), .left({trees[1771], lumberyards[1771]}), .right({trees[1773], lumberyards[1773]}), .bottom_left({trees[1821], lumberyards[1821]}), .bottom({trees[1822], lumberyards[1822]}), .bottom_right({trees[1823], lumberyards[1823]}), .init(2'b01), .state({trees[1772], lumberyards[1772]}));
acre acre_35_23 (.clk(clk), .en(en), .top_left({trees[1722], lumberyards[1722]}), .top({trees[1723], lumberyards[1723]}), .top_right({trees[1724], lumberyards[1724]}), .left({trees[1772], lumberyards[1772]}), .right({trees[1774], lumberyards[1774]}), .bottom_left({trees[1822], lumberyards[1822]}), .bottom({trees[1823], lumberyards[1823]}), .bottom_right({trees[1824], lumberyards[1824]}), .init(2'b00), .state({trees[1773], lumberyards[1773]}));
acre acre_35_24 (.clk(clk), .en(en), .top_left({trees[1723], lumberyards[1723]}), .top({trees[1724], lumberyards[1724]}), .top_right({trees[1725], lumberyards[1725]}), .left({trees[1773], lumberyards[1773]}), .right({trees[1775], lumberyards[1775]}), .bottom_left({trees[1823], lumberyards[1823]}), .bottom({trees[1824], lumberyards[1824]}), .bottom_right({trees[1825], lumberyards[1825]}), .init(2'b01), .state({trees[1774], lumberyards[1774]}));
acre acre_35_25 (.clk(clk), .en(en), .top_left({trees[1724], lumberyards[1724]}), .top({trees[1725], lumberyards[1725]}), .top_right({trees[1726], lumberyards[1726]}), .left({trees[1774], lumberyards[1774]}), .right({trees[1776], lumberyards[1776]}), .bottom_left({trees[1824], lumberyards[1824]}), .bottom({trees[1825], lumberyards[1825]}), .bottom_right({trees[1826], lumberyards[1826]}), .init(2'b10), .state({trees[1775], lumberyards[1775]}));
acre acre_35_26 (.clk(clk), .en(en), .top_left({trees[1725], lumberyards[1725]}), .top({trees[1726], lumberyards[1726]}), .top_right({trees[1727], lumberyards[1727]}), .left({trees[1775], lumberyards[1775]}), .right({trees[1777], lumberyards[1777]}), .bottom_left({trees[1825], lumberyards[1825]}), .bottom({trees[1826], lumberyards[1826]}), .bottom_right({trees[1827], lumberyards[1827]}), .init(2'b00), .state({trees[1776], lumberyards[1776]}));
acre acre_35_27 (.clk(clk), .en(en), .top_left({trees[1726], lumberyards[1726]}), .top({trees[1727], lumberyards[1727]}), .top_right({trees[1728], lumberyards[1728]}), .left({trees[1776], lumberyards[1776]}), .right({trees[1778], lumberyards[1778]}), .bottom_left({trees[1826], lumberyards[1826]}), .bottom({trees[1827], lumberyards[1827]}), .bottom_right({trees[1828], lumberyards[1828]}), .init(2'b00), .state({trees[1777], lumberyards[1777]}));
acre acre_35_28 (.clk(clk), .en(en), .top_left({trees[1727], lumberyards[1727]}), .top({trees[1728], lumberyards[1728]}), .top_right({trees[1729], lumberyards[1729]}), .left({trees[1777], lumberyards[1777]}), .right({trees[1779], lumberyards[1779]}), .bottom_left({trees[1827], lumberyards[1827]}), .bottom({trees[1828], lumberyards[1828]}), .bottom_right({trees[1829], lumberyards[1829]}), .init(2'b10), .state({trees[1778], lumberyards[1778]}));
acre acre_35_29 (.clk(clk), .en(en), .top_left({trees[1728], lumberyards[1728]}), .top({trees[1729], lumberyards[1729]}), .top_right({trees[1730], lumberyards[1730]}), .left({trees[1778], lumberyards[1778]}), .right({trees[1780], lumberyards[1780]}), .bottom_left({trees[1828], lumberyards[1828]}), .bottom({trees[1829], lumberyards[1829]}), .bottom_right({trees[1830], lumberyards[1830]}), .init(2'b01), .state({trees[1779], lumberyards[1779]}));
acre acre_35_30 (.clk(clk), .en(en), .top_left({trees[1729], lumberyards[1729]}), .top({trees[1730], lumberyards[1730]}), .top_right({trees[1731], lumberyards[1731]}), .left({trees[1779], lumberyards[1779]}), .right({trees[1781], lumberyards[1781]}), .bottom_left({trees[1829], lumberyards[1829]}), .bottom({trees[1830], lumberyards[1830]}), .bottom_right({trees[1831], lumberyards[1831]}), .init(2'b01), .state({trees[1780], lumberyards[1780]}));
acre acre_35_31 (.clk(clk), .en(en), .top_left({trees[1730], lumberyards[1730]}), .top({trees[1731], lumberyards[1731]}), .top_right({trees[1732], lumberyards[1732]}), .left({trees[1780], lumberyards[1780]}), .right({trees[1782], lumberyards[1782]}), .bottom_left({trees[1830], lumberyards[1830]}), .bottom({trees[1831], lumberyards[1831]}), .bottom_right({trees[1832], lumberyards[1832]}), .init(2'b10), .state({trees[1781], lumberyards[1781]}));
acre acre_35_32 (.clk(clk), .en(en), .top_left({trees[1731], lumberyards[1731]}), .top({trees[1732], lumberyards[1732]}), .top_right({trees[1733], lumberyards[1733]}), .left({trees[1781], lumberyards[1781]}), .right({trees[1783], lumberyards[1783]}), .bottom_left({trees[1831], lumberyards[1831]}), .bottom({trees[1832], lumberyards[1832]}), .bottom_right({trees[1833], lumberyards[1833]}), .init(2'b00), .state({trees[1782], lumberyards[1782]}));
acre acre_35_33 (.clk(clk), .en(en), .top_left({trees[1732], lumberyards[1732]}), .top({trees[1733], lumberyards[1733]}), .top_right({trees[1734], lumberyards[1734]}), .left({trees[1782], lumberyards[1782]}), .right({trees[1784], lumberyards[1784]}), .bottom_left({trees[1832], lumberyards[1832]}), .bottom({trees[1833], lumberyards[1833]}), .bottom_right({trees[1834], lumberyards[1834]}), .init(2'b01), .state({trees[1783], lumberyards[1783]}));
acre acre_35_34 (.clk(clk), .en(en), .top_left({trees[1733], lumberyards[1733]}), .top({trees[1734], lumberyards[1734]}), .top_right({trees[1735], lumberyards[1735]}), .left({trees[1783], lumberyards[1783]}), .right({trees[1785], lumberyards[1785]}), .bottom_left({trees[1833], lumberyards[1833]}), .bottom({trees[1834], lumberyards[1834]}), .bottom_right({trees[1835], lumberyards[1835]}), .init(2'b01), .state({trees[1784], lumberyards[1784]}));
acre acre_35_35 (.clk(clk), .en(en), .top_left({trees[1734], lumberyards[1734]}), .top({trees[1735], lumberyards[1735]}), .top_right({trees[1736], lumberyards[1736]}), .left({trees[1784], lumberyards[1784]}), .right({trees[1786], lumberyards[1786]}), .bottom_left({trees[1834], lumberyards[1834]}), .bottom({trees[1835], lumberyards[1835]}), .bottom_right({trees[1836], lumberyards[1836]}), .init(2'b00), .state({trees[1785], lumberyards[1785]}));
acre acre_35_36 (.clk(clk), .en(en), .top_left({trees[1735], lumberyards[1735]}), .top({trees[1736], lumberyards[1736]}), .top_right({trees[1737], lumberyards[1737]}), .left({trees[1785], lumberyards[1785]}), .right({trees[1787], lumberyards[1787]}), .bottom_left({trees[1835], lumberyards[1835]}), .bottom({trees[1836], lumberyards[1836]}), .bottom_right({trees[1837], lumberyards[1837]}), .init(2'b00), .state({trees[1786], lumberyards[1786]}));
acre acre_35_37 (.clk(clk), .en(en), .top_left({trees[1736], lumberyards[1736]}), .top({trees[1737], lumberyards[1737]}), .top_right({trees[1738], lumberyards[1738]}), .left({trees[1786], lumberyards[1786]}), .right({trees[1788], lumberyards[1788]}), .bottom_left({trees[1836], lumberyards[1836]}), .bottom({trees[1837], lumberyards[1837]}), .bottom_right({trees[1838], lumberyards[1838]}), .init(2'b00), .state({trees[1787], lumberyards[1787]}));
acre acre_35_38 (.clk(clk), .en(en), .top_left({trees[1737], lumberyards[1737]}), .top({trees[1738], lumberyards[1738]}), .top_right({trees[1739], lumberyards[1739]}), .left({trees[1787], lumberyards[1787]}), .right({trees[1789], lumberyards[1789]}), .bottom_left({trees[1837], lumberyards[1837]}), .bottom({trees[1838], lumberyards[1838]}), .bottom_right({trees[1839], lumberyards[1839]}), .init(2'b00), .state({trees[1788], lumberyards[1788]}));
acre acre_35_39 (.clk(clk), .en(en), .top_left({trees[1738], lumberyards[1738]}), .top({trees[1739], lumberyards[1739]}), .top_right({trees[1740], lumberyards[1740]}), .left({trees[1788], lumberyards[1788]}), .right({trees[1790], lumberyards[1790]}), .bottom_left({trees[1838], lumberyards[1838]}), .bottom({trees[1839], lumberyards[1839]}), .bottom_right({trees[1840], lumberyards[1840]}), .init(2'b01), .state({trees[1789], lumberyards[1789]}));
acre acre_35_40 (.clk(clk), .en(en), .top_left({trees[1739], lumberyards[1739]}), .top({trees[1740], lumberyards[1740]}), .top_right({trees[1741], lumberyards[1741]}), .left({trees[1789], lumberyards[1789]}), .right({trees[1791], lumberyards[1791]}), .bottom_left({trees[1839], lumberyards[1839]}), .bottom({trees[1840], lumberyards[1840]}), .bottom_right({trees[1841], lumberyards[1841]}), .init(2'b00), .state({trees[1790], lumberyards[1790]}));
acre acre_35_41 (.clk(clk), .en(en), .top_left({trees[1740], lumberyards[1740]}), .top({trees[1741], lumberyards[1741]}), .top_right({trees[1742], lumberyards[1742]}), .left({trees[1790], lumberyards[1790]}), .right({trees[1792], lumberyards[1792]}), .bottom_left({trees[1840], lumberyards[1840]}), .bottom({trees[1841], lumberyards[1841]}), .bottom_right({trees[1842], lumberyards[1842]}), .init(2'b01), .state({trees[1791], lumberyards[1791]}));
acre acre_35_42 (.clk(clk), .en(en), .top_left({trees[1741], lumberyards[1741]}), .top({trees[1742], lumberyards[1742]}), .top_right({trees[1743], lumberyards[1743]}), .left({trees[1791], lumberyards[1791]}), .right({trees[1793], lumberyards[1793]}), .bottom_left({trees[1841], lumberyards[1841]}), .bottom({trees[1842], lumberyards[1842]}), .bottom_right({trees[1843], lumberyards[1843]}), .init(2'b01), .state({trees[1792], lumberyards[1792]}));
acre acre_35_43 (.clk(clk), .en(en), .top_left({trees[1742], lumberyards[1742]}), .top({trees[1743], lumberyards[1743]}), .top_right({trees[1744], lumberyards[1744]}), .left({trees[1792], lumberyards[1792]}), .right({trees[1794], lumberyards[1794]}), .bottom_left({trees[1842], lumberyards[1842]}), .bottom({trees[1843], lumberyards[1843]}), .bottom_right({trees[1844], lumberyards[1844]}), .init(2'b10), .state({trees[1793], lumberyards[1793]}));
acre acre_35_44 (.clk(clk), .en(en), .top_left({trees[1743], lumberyards[1743]}), .top({trees[1744], lumberyards[1744]}), .top_right({trees[1745], lumberyards[1745]}), .left({trees[1793], lumberyards[1793]}), .right({trees[1795], lumberyards[1795]}), .bottom_left({trees[1843], lumberyards[1843]}), .bottom({trees[1844], lumberyards[1844]}), .bottom_right({trees[1845], lumberyards[1845]}), .init(2'b00), .state({trees[1794], lumberyards[1794]}));
acre acre_35_45 (.clk(clk), .en(en), .top_left({trees[1744], lumberyards[1744]}), .top({trees[1745], lumberyards[1745]}), .top_right({trees[1746], lumberyards[1746]}), .left({trees[1794], lumberyards[1794]}), .right({trees[1796], lumberyards[1796]}), .bottom_left({trees[1844], lumberyards[1844]}), .bottom({trees[1845], lumberyards[1845]}), .bottom_right({trees[1846], lumberyards[1846]}), .init(2'b00), .state({trees[1795], lumberyards[1795]}));
acre acre_35_46 (.clk(clk), .en(en), .top_left({trees[1745], lumberyards[1745]}), .top({trees[1746], lumberyards[1746]}), .top_right({trees[1747], lumberyards[1747]}), .left({trees[1795], lumberyards[1795]}), .right({trees[1797], lumberyards[1797]}), .bottom_left({trees[1845], lumberyards[1845]}), .bottom({trees[1846], lumberyards[1846]}), .bottom_right({trees[1847], lumberyards[1847]}), .init(2'b00), .state({trees[1796], lumberyards[1796]}));
acre acre_35_47 (.clk(clk), .en(en), .top_left({trees[1746], lumberyards[1746]}), .top({trees[1747], lumberyards[1747]}), .top_right({trees[1748], lumberyards[1748]}), .left({trees[1796], lumberyards[1796]}), .right({trees[1798], lumberyards[1798]}), .bottom_left({trees[1846], lumberyards[1846]}), .bottom({trees[1847], lumberyards[1847]}), .bottom_right({trees[1848], lumberyards[1848]}), .init(2'b00), .state({trees[1797], lumberyards[1797]}));
acre acre_35_48 (.clk(clk), .en(en), .top_left({trees[1747], lumberyards[1747]}), .top({trees[1748], lumberyards[1748]}), .top_right({trees[1749], lumberyards[1749]}), .left({trees[1797], lumberyards[1797]}), .right({trees[1799], lumberyards[1799]}), .bottom_left({trees[1847], lumberyards[1847]}), .bottom({trees[1848], lumberyards[1848]}), .bottom_right({trees[1849], lumberyards[1849]}), .init(2'b10), .state({trees[1798], lumberyards[1798]}));
acre acre_35_49 (.clk(clk), .en(en), .top_left({trees[1748], lumberyards[1748]}), .top({trees[1749], lumberyards[1749]}), .top_right(2'b0), .left({trees[1798], lumberyards[1798]}), .right(2'b0), .bottom_left({trees[1848], lumberyards[1848]}), .bottom({trees[1849], lumberyards[1849]}), .bottom_right(2'b0), .init(2'b00), .state({trees[1799], lumberyards[1799]}));
acre acre_36_0 (.clk(clk), .en(en), .top_left(2'b0), .top({trees[1750], lumberyards[1750]}), .top_right({trees[1751], lumberyards[1751]}), .left(2'b0), .right({trees[1801], lumberyards[1801]}), .bottom_left(2'b0), .bottom({trees[1850], lumberyards[1850]}), .bottom_right({trees[1851], lumberyards[1851]}), .init(2'b00), .state({trees[1800], lumberyards[1800]}));
acre acre_36_1 (.clk(clk), .en(en), .top_left({trees[1750], lumberyards[1750]}), .top({trees[1751], lumberyards[1751]}), .top_right({trees[1752], lumberyards[1752]}), .left({trees[1800], lumberyards[1800]}), .right({trees[1802], lumberyards[1802]}), .bottom_left({trees[1850], lumberyards[1850]}), .bottom({trees[1851], lumberyards[1851]}), .bottom_right({trees[1852], lumberyards[1852]}), .init(2'b10), .state({trees[1801], lumberyards[1801]}));
acre acre_36_2 (.clk(clk), .en(en), .top_left({trees[1751], lumberyards[1751]}), .top({trees[1752], lumberyards[1752]}), .top_right({trees[1753], lumberyards[1753]}), .left({trees[1801], lumberyards[1801]}), .right({trees[1803], lumberyards[1803]}), .bottom_left({trees[1851], lumberyards[1851]}), .bottom({trees[1852], lumberyards[1852]}), .bottom_right({trees[1853], lumberyards[1853]}), .init(2'b10), .state({trees[1802], lumberyards[1802]}));
acre acre_36_3 (.clk(clk), .en(en), .top_left({trees[1752], lumberyards[1752]}), .top({trees[1753], lumberyards[1753]}), .top_right({trees[1754], lumberyards[1754]}), .left({trees[1802], lumberyards[1802]}), .right({trees[1804], lumberyards[1804]}), .bottom_left({trees[1852], lumberyards[1852]}), .bottom({trees[1853], lumberyards[1853]}), .bottom_right({trees[1854], lumberyards[1854]}), .init(2'b00), .state({trees[1803], lumberyards[1803]}));
acre acre_36_4 (.clk(clk), .en(en), .top_left({trees[1753], lumberyards[1753]}), .top({trees[1754], lumberyards[1754]}), .top_right({trees[1755], lumberyards[1755]}), .left({trees[1803], lumberyards[1803]}), .right({trees[1805], lumberyards[1805]}), .bottom_left({trees[1853], lumberyards[1853]}), .bottom({trees[1854], lumberyards[1854]}), .bottom_right({trees[1855], lumberyards[1855]}), .init(2'b00), .state({trees[1804], lumberyards[1804]}));
acre acre_36_5 (.clk(clk), .en(en), .top_left({trees[1754], lumberyards[1754]}), .top({trees[1755], lumberyards[1755]}), .top_right({trees[1756], lumberyards[1756]}), .left({trees[1804], lumberyards[1804]}), .right({trees[1806], lumberyards[1806]}), .bottom_left({trees[1854], lumberyards[1854]}), .bottom({trees[1855], lumberyards[1855]}), .bottom_right({trees[1856], lumberyards[1856]}), .init(2'b00), .state({trees[1805], lumberyards[1805]}));
acre acre_36_6 (.clk(clk), .en(en), .top_left({trees[1755], lumberyards[1755]}), .top({trees[1756], lumberyards[1756]}), .top_right({trees[1757], lumberyards[1757]}), .left({trees[1805], lumberyards[1805]}), .right({trees[1807], lumberyards[1807]}), .bottom_left({trees[1855], lumberyards[1855]}), .bottom({trees[1856], lumberyards[1856]}), .bottom_right({trees[1857], lumberyards[1857]}), .init(2'b10), .state({trees[1806], lumberyards[1806]}));
acre acre_36_7 (.clk(clk), .en(en), .top_left({trees[1756], lumberyards[1756]}), .top({trees[1757], lumberyards[1757]}), .top_right({trees[1758], lumberyards[1758]}), .left({trees[1806], lumberyards[1806]}), .right({trees[1808], lumberyards[1808]}), .bottom_left({trees[1856], lumberyards[1856]}), .bottom({trees[1857], lumberyards[1857]}), .bottom_right({trees[1858], lumberyards[1858]}), .init(2'b10), .state({trees[1807], lumberyards[1807]}));
acre acre_36_8 (.clk(clk), .en(en), .top_left({trees[1757], lumberyards[1757]}), .top({trees[1758], lumberyards[1758]}), .top_right({trees[1759], lumberyards[1759]}), .left({trees[1807], lumberyards[1807]}), .right({trees[1809], lumberyards[1809]}), .bottom_left({trees[1857], lumberyards[1857]}), .bottom({trees[1858], lumberyards[1858]}), .bottom_right({trees[1859], lumberyards[1859]}), .init(2'b00), .state({trees[1808], lumberyards[1808]}));
acre acre_36_9 (.clk(clk), .en(en), .top_left({trees[1758], lumberyards[1758]}), .top({trees[1759], lumberyards[1759]}), .top_right({trees[1760], lumberyards[1760]}), .left({trees[1808], lumberyards[1808]}), .right({trees[1810], lumberyards[1810]}), .bottom_left({trees[1858], lumberyards[1858]}), .bottom({trees[1859], lumberyards[1859]}), .bottom_right({trees[1860], lumberyards[1860]}), .init(2'b10), .state({trees[1809], lumberyards[1809]}));
acre acre_36_10 (.clk(clk), .en(en), .top_left({trees[1759], lumberyards[1759]}), .top({trees[1760], lumberyards[1760]}), .top_right({trees[1761], lumberyards[1761]}), .left({trees[1809], lumberyards[1809]}), .right({trees[1811], lumberyards[1811]}), .bottom_left({trees[1859], lumberyards[1859]}), .bottom({trees[1860], lumberyards[1860]}), .bottom_right({trees[1861], lumberyards[1861]}), .init(2'b00), .state({trees[1810], lumberyards[1810]}));
acre acre_36_11 (.clk(clk), .en(en), .top_left({trees[1760], lumberyards[1760]}), .top({trees[1761], lumberyards[1761]}), .top_right({trees[1762], lumberyards[1762]}), .left({trees[1810], lumberyards[1810]}), .right({trees[1812], lumberyards[1812]}), .bottom_left({trees[1860], lumberyards[1860]}), .bottom({trees[1861], lumberyards[1861]}), .bottom_right({trees[1862], lumberyards[1862]}), .init(2'b00), .state({trees[1811], lumberyards[1811]}));
acre acre_36_12 (.clk(clk), .en(en), .top_left({trees[1761], lumberyards[1761]}), .top({trees[1762], lumberyards[1762]}), .top_right({trees[1763], lumberyards[1763]}), .left({trees[1811], lumberyards[1811]}), .right({trees[1813], lumberyards[1813]}), .bottom_left({trees[1861], lumberyards[1861]}), .bottom({trees[1862], lumberyards[1862]}), .bottom_right({trees[1863], lumberyards[1863]}), .init(2'b01), .state({trees[1812], lumberyards[1812]}));
acre acre_36_13 (.clk(clk), .en(en), .top_left({trees[1762], lumberyards[1762]}), .top({trees[1763], lumberyards[1763]}), .top_right({trees[1764], lumberyards[1764]}), .left({trees[1812], lumberyards[1812]}), .right({trees[1814], lumberyards[1814]}), .bottom_left({trees[1862], lumberyards[1862]}), .bottom({trees[1863], lumberyards[1863]}), .bottom_right({trees[1864], lumberyards[1864]}), .init(2'b00), .state({trees[1813], lumberyards[1813]}));
acre acre_36_14 (.clk(clk), .en(en), .top_left({trees[1763], lumberyards[1763]}), .top({trees[1764], lumberyards[1764]}), .top_right({trees[1765], lumberyards[1765]}), .left({trees[1813], lumberyards[1813]}), .right({trees[1815], lumberyards[1815]}), .bottom_left({trees[1863], lumberyards[1863]}), .bottom({trees[1864], lumberyards[1864]}), .bottom_right({trees[1865], lumberyards[1865]}), .init(2'b00), .state({trees[1814], lumberyards[1814]}));
acre acre_36_15 (.clk(clk), .en(en), .top_left({trees[1764], lumberyards[1764]}), .top({trees[1765], lumberyards[1765]}), .top_right({trees[1766], lumberyards[1766]}), .left({trees[1814], lumberyards[1814]}), .right({trees[1816], lumberyards[1816]}), .bottom_left({trees[1864], lumberyards[1864]}), .bottom({trees[1865], lumberyards[1865]}), .bottom_right({trees[1866], lumberyards[1866]}), .init(2'b00), .state({trees[1815], lumberyards[1815]}));
acre acre_36_16 (.clk(clk), .en(en), .top_left({trees[1765], lumberyards[1765]}), .top({trees[1766], lumberyards[1766]}), .top_right({trees[1767], lumberyards[1767]}), .left({trees[1815], lumberyards[1815]}), .right({trees[1817], lumberyards[1817]}), .bottom_left({trees[1865], lumberyards[1865]}), .bottom({trees[1866], lumberyards[1866]}), .bottom_right({trees[1867], lumberyards[1867]}), .init(2'b00), .state({trees[1816], lumberyards[1816]}));
acre acre_36_17 (.clk(clk), .en(en), .top_left({trees[1766], lumberyards[1766]}), .top({trees[1767], lumberyards[1767]}), .top_right({trees[1768], lumberyards[1768]}), .left({trees[1816], lumberyards[1816]}), .right({trees[1818], lumberyards[1818]}), .bottom_left({trees[1866], lumberyards[1866]}), .bottom({trees[1867], lumberyards[1867]}), .bottom_right({trees[1868], lumberyards[1868]}), .init(2'b10), .state({trees[1817], lumberyards[1817]}));
acre acre_36_18 (.clk(clk), .en(en), .top_left({trees[1767], lumberyards[1767]}), .top({trees[1768], lumberyards[1768]}), .top_right({trees[1769], lumberyards[1769]}), .left({trees[1817], lumberyards[1817]}), .right({trees[1819], lumberyards[1819]}), .bottom_left({trees[1867], lumberyards[1867]}), .bottom({trees[1868], lumberyards[1868]}), .bottom_right({trees[1869], lumberyards[1869]}), .init(2'b10), .state({trees[1818], lumberyards[1818]}));
acre acre_36_19 (.clk(clk), .en(en), .top_left({trees[1768], lumberyards[1768]}), .top({trees[1769], lumberyards[1769]}), .top_right({trees[1770], lumberyards[1770]}), .left({trees[1818], lumberyards[1818]}), .right({trees[1820], lumberyards[1820]}), .bottom_left({trees[1868], lumberyards[1868]}), .bottom({trees[1869], lumberyards[1869]}), .bottom_right({trees[1870], lumberyards[1870]}), .init(2'b00), .state({trees[1819], lumberyards[1819]}));
acre acre_36_20 (.clk(clk), .en(en), .top_left({trees[1769], lumberyards[1769]}), .top({trees[1770], lumberyards[1770]}), .top_right({trees[1771], lumberyards[1771]}), .left({trees[1819], lumberyards[1819]}), .right({trees[1821], lumberyards[1821]}), .bottom_left({trees[1869], lumberyards[1869]}), .bottom({trees[1870], lumberyards[1870]}), .bottom_right({trees[1871], lumberyards[1871]}), .init(2'b00), .state({trees[1820], lumberyards[1820]}));
acre acre_36_21 (.clk(clk), .en(en), .top_left({trees[1770], lumberyards[1770]}), .top({trees[1771], lumberyards[1771]}), .top_right({trees[1772], lumberyards[1772]}), .left({trees[1820], lumberyards[1820]}), .right({trees[1822], lumberyards[1822]}), .bottom_left({trees[1870], lumberyards[1870]}), .bottom({trees[1871], lumberyards[1871]}), .bottom_right({trees[1872], lumberyards[1872]}), .init(2'b10), .state({trees[1821], lumberyards[1821]}));
acre acre_36_22 (.clk(clk), .en(en), .top_left({trees[1771], lumberyards[1771]}), .top({trees[1772], lumberyards[1772]}), .top_right({trees[1773], lumberyards[1773]}), .left({trees[1821], lumberyards[1821]}), .right({trees[1823], lumberyards[1823]}), .bottom_left({trees[1871], lumberyards[1871]}), .bottom({trees[1872], lumberyards[1872]}), .bottom_right({trees[1873], lumberyards[1873]}), .init(2'b01), .state({trees[1822], lumberyards[1822]}));
acre acre_36_23 (.clk(clk), .en(en), .top_left({trees[1772], lumberyards[1772]}), .top({trees[1773], lumberyards[1773]}), .top_right({trees[1774], lumberyards[1774]}), .left({trees[1822], lumberyards[1822]}), .right({trees[1824], lumberyards[1824]}), .bottom_left({trees[1872], lumberyards[1872]}), .bottom({trees[1873], lumberyards[1873]}), .bottom_right({trees[1874], lumberyards[1874]}), .init(2'b00), .state({trees[1823], lumberyards[1823]}));
acre acre_36_24 (.clk(clk), .en(en), .top_left({trees[1773], lumberyards[1773]}), .top({trees[1774], lumberyards[1774]}), .top_right({trees[1775], lumberyards[1775]}), .left({trees[1823], lumberyards[1823]}), .right({trees[1825], lumberyards[1825]}), .bottom_left({trees[1873], lumberyards[1873]}), .bottom({trees[1874], lumberyards[1874]}), .bottom_right({trees[1875], lumberyards[1875]}), .init(2'b00), .state({trees[1824], lumberyards[1824]}));
acre acre_36_25 (.clk(clk), .en(en), .top_left({trees[1774], lumberyards[1774]}), .top({trees[1775], lumberyards[1775]}), .top_right({trees[1776], lumberyards[1776]}), .left({trees[1824], lumberyards[1824]}), .right({trees[1826], lumberyards[1826]}), .bottom_left({trees[1874], lumberyards[1874]}), .bottom({trees[1875], lumberyards[1875]}), .bottom_right({trees[1876], lumberyards[1876]}), .init(2'b00), .state({trees[1825], lumberyards[1825]}));
acre acre_36_26 (.clk(clk), .en(en), .top_left({trees[1775], lumberyards[1775]}), .top({trees[1776], lumberyards[1776]}), .top_right({trees[1777], lumberyards[1777]}), .left({trees[1825], lumberyards[1825]}), .right({trees[1827], lumberyards[1827]}), .bottom_left({trees[1875], lumberyards[1875]}), .bottom({trees[1876], lumberyards[1876]}), .bottom_right({trees[1877], lumberyards[1877]}), .init(2'b10), .state({trees[1826], lumberyards[1826]}));
acre acre_36_27 (.clk(clk), .en(en), .top_left({trees[1776], lumberyards[1776]}), .top({trees[1777], lumberyards[1777]}), .top_right({trees[1778], lumberyards[1778]}), .left({trees[1826], lumberyards[1826]}), .right({trees[1828], lumberyards[1828]}), .bottom_left({trees[1876], lumberyards[1876]}), .bottom({trees[1877], lumberyards[1877]}), .bottom_right({trees[1878], lumberyards[1878]}), .init(2'b01), .state({trees[1827], lumberyards[1827]}));
acre acre_36_28 (.clk(clk), .en(en), .top_left({trees[1777], lumberyards[1777]}), .top({trees[1778], lumberyards[1778]}), .top_right({trees[1779], lumberyards[1779]}), .left({trees[1827], lumberyards[1827]}), .right({trees[1829], lumberyards[1829]}), .bottom_left({trees[1877], lumberyards[1877]}), .bottom({trees[1878], lumberyards[1878]}), .bottom_right({trees[1879], lumberyards[1879]}), .init(2'b01), .state({trees[1828], lumberyards[1828]}));
acre acre_36_29 (.clk(clk), .en(en), .top_left({trees[1778], lumberyards[1778]}), .top({trees[1779], lumberyards[1779]}), .top_right({trees[1780], lumberyards[1780]}), .left({trees[1828], lumberyards[1828]}), .right({trees[1830], lumberyards[1830]}), .bottom_left({trees[1878], lumberyards[1878]}), .bottom({trees[1879], lumberyards[1879]}), .bottom_right({trees[1880], lumberyards[1880]}), .init(2'b01), .state({trees[1829], lumberyards[1829]}));
acre acre_36_30 (.clk(clk), .en(en), .top_left({trees[1779], lumberyards[1779]}), .top({trees[1780], lumberyards[1780]}), .top_right({trees[1781], lumberyards[1781]}), .left({trees[1829], lumberyards[1829]}), .right({trees[1831], lumberyards[1831]}), .bottom_left({trees[1879], lumberyards[1879]}), .bottom({trees[1880], lumberyards[1880]}), .bottom_right({trees[1881], lumberyards[1881]}), .init(2'b00), .state({trees[1830], lumberyards[1830]}));
acre acre_36_31 (.clk(clk), .en(en), .top_left({trees[1780], lumberyards[1780]}), .top({trees[1781], lumberyards[1781]}), .top_right({trees[1782], lumberyards[1782]}), .left({trees[1830], lumberyards[1830]}), .right({trees[1832], lumberyards[1832]}), .bottom_left({trees[1880], lumberyards[1880]}), .bottom({trees[1881], lumberyards[1881]}), .bottom_right({trees[1882], lumberyards[1882]}), .init(2'b00), .state({trees[1831], lumberyards[1831]}));
acre acre_36_32 (.clk(clk), .en(en), .top_left({trees[1781], lumberyards[1781]}), .top({trees[1782], lumberyards[1782]}), .top_right({trees[1783], lumberyards[1783]}), .left({trees[1831], lumberyards[1831]}), .right({trees[1833], lumberyards[1833]}), .bottom_left({trees[1881], lumberyards[1881]}), .bottom({trees[1882], lumberyards[1882]}), .bottom_right({trees[1883], lumberyards[1883]}), .init(2'b01), .state({trees[1832], lumberyards[1832]}));
acre acre_36_33 (.clk(clk), .en(en), .top_left({trees[1782], lumberyards[1782]}), .top({trees[1783], lumberyards[1783]}), .top_right({trees[1784], lumberyards[1784]}), .left({trees[1832], lumberyards[1832]}), .right({trees[1834], lumberyards[1834]}), .bottom_left({trees[1882], lumberyards[1882]}), .bottom({trees[1883], lumberyards[1883]}), .bottom_right({trees[1884], lumberyards[1884]}), .init(2'b00), .state({trees[1833], lumberyards[1833]}));
acre acre_36_34 (.clk(clk), .en(en), .top_left({trees[1783], lumberyards[1783]}), .top({trees[1784], lumberyards[1784]}), .top_right({trees[1785], lumberyards[1785]}), .left({trees[1833], lumberyards[1833]}), .right({trees[1835], lumberyards[1835]}), .bottom_left({trees[1883], lumberyards[1883]}), .bottom({trees[1884], lumberyards[1884]}), .bottom_right({trees[1885], lumberyards[1885]}), .init(2'b00), .state({trees[1834], lumberyards[1834]}));
acre acre_36_35 (.clk(clk), .en(en), .top_left({trees[1784], lumberyards[1784]}), .top({trees[1785], lumberyards[1785]}), .top_right({trees[1786], lumberyards[1786]}), .left({trees[1834], lumberyards[1834]}), .right({trees[1836], lumberyards[1836]}), .bottom_left({trees[1884], lumberyards[1884]}), .bottom({trees[1885], lumberyards[1885]}), .bottom_right({trees[1886], lumberyards[1886]}), .init(2'b00), .state({trees[1835], lumberyards[1835]}));
acre acre_36_36 (.clk(clk), .en(en), .top_left({trees[1785], lumberyards[1785]}), .top({trees[1786], lumberyards[1786]}), .top_right({trees[1787], lumberyards[1787]}), .left({trees[1835], lumberyards[1835]}), .right({trees[1837], lumberyards[1837]}), .bottom_left({trees[1885], lumberyards[1885]}), .bottom({trees[1886], lumberyards[1886]}), .bottom_right({trees[1887], lumberyards[1887]}), .init(2'b00), .state({trees[1836], lumberyards[1836]}));
acre acre_36_37 (.clk(clk), .en(en), .top_left({trees[1786], lumberyards[1786]}), .top({trees[1787], lumberyards[1787]}), .top_right({trees[1788], lumberyards[1788]}), .left({trees[1836], lumberyards[1836]}), .right({trees[1838], lumberyards[1838]}), .bottom_left({trees[1886], lumberyards[1886]}), .bottom({trees[1887], lumberyards[1887]}), .bottom_right({trees[1888], lumberyards[1888]}), .init(2'b01), .state({trees[1837], lumberyards[1837]}));
acre acre_36_38 (.clk(clk), .en(en), .top_left({trees[1787], lumberyards[1787]}), .top({trees[1788], lumberyards[1788]}), .top_right({trees[1789], lumberyards[1789]}), .left({trees[1837], lumberyards[1837]}), .right({trees[1839], lumberyards[1839]}), .bottom_left({trees[1887], lumberyards[1887]}), .bottom({trees[1888], lumberyards[1888]}), .bottom_right({trees[1889], lumberyards[1889]}), .init(2'b00), .state({trees[1838], lumberyards[1838]}));
acre acre_36_39 (.clk(clk), .en(en), .top_left({trees[1788], lumberyards[1788]}), .top({trees[1789], lumberyards[1789]}), .top_right({trees[1790], lumberyards[1790]}), .left({trees[1838], lumberyards[1838]}), .right({trees[1840], lumberyards[1840]}), .bottom_left({trees[1888], lumberyards[1888]}), .bottom({trees[1889], lumberyards[1889]}), .bottom_right({trees[1890], lumberyards[1890]}), .init(2'b01), .state({trees[1839], lumberyards[1839]}));
acre acre_36_40 (.clk(clk), .en(en), .top_left({trees[1789], lumberyards[1789]}), .top({trees[1790], lumberyards[1790]}), .top_right({trees[1791], lumberyards[1791]}), .left({trees[1839], lumberyards[1839]}), .right({trees[1841], lumberyards[1841]}), .bottom_left({trees[1889], lumberyards[1889]}), .bottom({trees[1890], lumberyards[1890]}), .bottom_right({trees[1891], lumberyards[1891]}), .init(2'b00), .state({trees[1840], lumberyards[1840]}));
acre acre_36_41 (.clk(clk), .en(en), .top_left({trees[1790], lumberyards[1790]}), .top({trees[1791], lumberyards[1791]}), .top_right({trees[1792], lumberyards[1792]}), .left({trees[1840], lumberyards[1840]}), .right({trees[1842], lumberyards[1842]}), .bottom_left({trees[1890], lumberyards[1890]}), .bottom({trees[1891], lumberyards[1891]}), .bottom_right({trees[1892], lumberyards[1892]}), .init(2'b00), .state({trees[1841], lumberyards[1841]}));
acre acre_36_42 (.clk(clk), .en(en), .top_left({trees[1791], lumberyards[1791]}), .top({trees[1792], lumberyards[1792]}), .top_right({trees[1793], lumberyards[1793]}), .left({trees[1841], lumberyards[1841]}), .right({trees[1843], lumberyards[1843]}), .bottom_left({trees[1891], lumberyards[1891]}), .bottom({trees[1892], lumberyards[1892]}), .bottom_right({trees[1893], lumberyards[1893]}), .init(2'b00), .state({trees[1842], lumberyards[1842]}));
acre acre_36_43 (.clk(clk), .en(en), .top_left({trees[1792], lumberyards[1792]}), .top({trees[1793], lumberyards[1793]}), .top_right({trees[1794], lumberyards[1794]}), .left({trees[1842], lumberyards[1842]}), .right({trees[1844], lumberyards[1844]}), .bottom_left({trees[1892], lumberyards[1892]}), .bottom({trees[1893], lumberyards[1893]}), .bottom_right({trees[1894], lumberyards[1894]}), .init(2'b00), .state({trees[1843], lumberyards[1843]}));
acre acre_36_44 (.clk(clk), .en(en), .top_left({trees[1793], lumberyards[1793]}), .top({trees[1794], lumberyards[1794]}), .top_right({trees[1795], lumberyards[1795]}), .left({trees[1843], lumberyards[1843]}), .right({trees[1845], lumberyards[1845]}), .bottom_left({trees[1893], lumberyards[1893]}), .bottom({trees[1894], lumberyards[1894]}), .bottom_right({trees[1895], lumberyards[1895]}), .init(2'b00), .state({trees[1844], lumberyards[1844]}));
acre acre_36_45 (.clk(clk), .en(en), .top_left({trees[1794], lumberyards[1794]}), .top({trees[1795], lumberyards[1795]}), .top_right({trees[1796], lumberyards[1796]}), .left({trees[1844], lumberyards[1844]}), .right({trees[1846], lumberyards[1846]}), .bottom_left({trees[1894], lumberyards[1894]}), .bottom({trees[1895], lumberyards[1895]}), .bottom_right({trees[1896], lumberyards[1896]}), .init(2'b00), .state({trees[1845], lumberyards[1845]}));
acre acre_36_46 (.clk(clk), .en(en), .top_left({trees[1795], lumberyards[1795]}), .top({trees[1796], lumberyards[1796]}), .top_right({trees[1797], lumberyards[1797]}), .left({trees[1845], lumberyards[1845]}), .right({trees[1847], lumberyards[1847]}), .bottom_left({trees[1895], lumberyards[1895]}), .bottom({trees[1896], lumberyards[1896]}), .bottom_right({trees[1897], lumberyards[1897]}), .init(2'b00), .state({trees[1846], lumberyards[1846]}));
acre acre_36_47 (.clk(clk), .en(en), .top_left({trees[1796], lumberyards[1796]}), .top({trees[1797], lumberyards[1797]}), .top_right({trees[1798], lumberyards[1798]}), .left({trees[1846], lumberyards[1846]}), .right({trees[1848], lumberyards[1848]}), .bottom_left({trees[1896], lumberyards[1896]}), .bottom({trees[1897], lumberyards[1897]}), .bottom_right({trees[1898], lumberyards[1898]}), .init(2'b10), .state({trees[1847], lumberyards[1847]}));
acre acre_36_48 (.clk(clk), .en(en), .top_left({trees[1797], lumberyards[1797]}), .top({trees[1798], lumberyards[1798]}), .top_right({trees[1799], lumberyards[1799]}), .left({trees[1847], lumberyards[1847]}), .right({trees[1849], lumberyards[1849]}), .bottom_left({trees[1897], lumberyards[1897]}), .bottom({trees[1898], lumberyards[1898]}), .bottom_right({trees[1899], lumberyards[1899]}), .init(2'b01), .state({trees[1848], lumberyards[1848]}));
acre acre_36_49 (.clk(clk), .en(en), .top_left({trees[1798], lumberyards[1798]}), .top({trees[1799], lumberyards[1799]}), .top_right(2'b0), .left({trees[1848], lumberyards[1848]}), .right(2'b0), .bottom_left({trees[1898], lumberyards[1898]}), .bottom({trees[1899], lumberyards[1899]}), .bottom_right(2'b0), .init(2'b00), .state({trees[1849], lumberyards[1849]}));
acre acre_37_0 (.clk(clk), .en(en), .top_left(2'b0), .top({trees[1800], lumberyards[1800]}), .top_right({trees[1801], lumberyards[1801]}), .left(2'b0), .right({trees[1851], lumberyards[1851]}), .bottom_left(2'b0), .bottom({trees[1900], lumberyards[1900]}), .bottom_right({trees[1901], lumberyards[1901]}), .init(2'b00), .state({trees[1850], lumberyards[1850]}));
acre acre_37_1 (.clk(clk), .en(en), .top_left({trees[1800], lumberyards[1800]}), .top({trees[1801], lumberyards[1801]}), .top_right({trees[1802], lumberyards[1802]}), .left({trees[1850], lumberyards[1850]}), .right({trees[1852], lumberyards[1852]}), .bottom_left({trees[1900], lumberyards[1900]}), .bottom({trees[1901], lumberyards[1901]}), .bottom_right({trees[1902], lumberyards[1902]}), .init(2'b10), .state({trees[1851], lumberyards[1851]}));
acre acre_37_2 (.clk(clk), .en(en), .top_left({trees[1801], lumberyards[1801]}), .top({trees[1802], lumberyards[1802]}), .top_right({trees[1803], lumberyards[1803]}), .left({trees[1851], lumberyards[1851]}), .right({trees[1853], lumberyards[1853]}), .bottom_left({trees[1901], lumberyards[1901]}), .bottom({trees[1902], lumberyards[1902]}), .bottom_right({trees[1903], lumberyards[1903]}), .init(2'b10), .state({trees[1852], lumberyards[1852]}));
acre acre_37_3 (.clk(clk), .en(en), .top_left({trees[1802], lumberyards[1802]}), .top({trees[1803], lumberyards[1803]}), .top_right({trees[1804], lumberyards[1804]}), .left({trees[1852], lumberyards[1852]}), .right({trees[1854], lumberyards[1854]}), .bottom_left({trees[1902], lumberyards[1902]}), .bottom({trees[1903], lumberyards[1903]}), .bottom_right({trees[1904], lumberyards[1904]}), .init(2'b01), .state({trees[1853], lumberyards[1853]}));
acre acre_37_4 (.clk(clk), .en(en), .top_left({trees[1803], lumberyards[1803]}), .top({trees[1804], lumberyards[1804]}), .top_right({trees[1805], lumberyards[1805]}), .left({trees[1853], lumberyards[1853]}), .right({trees[1855], lumberyards[1855]}), .bottom_left({trees[1903], lumberyards[1903]}), .bottom({trees[1904], lumberyards[1904]}), .bottom_right({trees[1905], lumberyards[1905]}), .init(2'b00), .state({trees[1854], lumberyards[1854]}));
acre acre_37_5 (.clk(clk), .en(en), .top_left({trees[1804], lumberyards[1804]}), .top({trees[1805], lumberyards[1805]}), .top_right({trees[1806], lumberyards[1806]}), .left({trees[1854], lumberyards[1854]}), .right({trees[1856], lumberyards[1856]}), .bottom_left({trees[1904], lumberyards[1904]}), .bottom({trees[1905], lumberyards[1905]}), .bottom_right({trees[1906], lumberyards[1906]}), .init(2'b10), .state({trees[1855], lumberyards[1855]}));
acre acre_37_6 (.clk(clk), .en(en), .top_left({trees[1805], lumberyards[1805]}), .top({trees[1806], lumberyards[1806]}), .top_right({trees[1807], lumberyards[1807]}), .left({trees[1855], lumberyards[1855]}), .right({trees[1857], lumberyards[1857]}), .bottom_left({trees[1905], lumberyards[1905]}), .bottom({trees[1906], lumberyards[1906]}), .bottom_right({trees[1907], lumberyards[1907]}), .init(2'b00), .state({trees[1856], lumberyards[1856]}));
acre acre_37_7 (.clk(clk), .en(en), .top_left({trees[1806], lumberyards[1806]}), .top({trees[1807], lumberyards[1807]}), .top_right({trees[1808], lumberyards[1808]}), .left({trees[1856], lumberyards[1856]}), .right({trees[1858], lumberyards[1858]}), .bottom_left({trees[1906], lumberyards[1906]}), .bottom({trees[1907], lumberyards[1907]}), .bottom_right({trees[1908], lumberyards[1908]}), .init(2'b00), .state({trees[1857], lumberyards[1857]}));
acre acre_37_8 (.clk(clk), .en(en), .top_left({trees[1807], lumberyards[1807]}), .top({trees[1808], lumberyards[1808]}), .top_right({trees[1809], lumberyards[1809]}), .left({trees[1857], lumberyards[1857]}), .right({trees[1859], lumberyards[1859]}), .bottom_left({trees[1907], lumberyards[1907]}), .bottom({trees[1908], lumberyards[1908]}), .bottom_right({trees[1909], lumberyards[1909]}), .init(2'b00), .state({trees[1858], lumberyards[1858]}));
acre acre_37_9 (.clk(clk), .en(en), .top_left({trees[1808], lumberyards[1808]}), .top({trees[1809], lumberyards[1809]}), .top_right({trees[1810], lumberyards[1810]}), .left({trees[1858], lumberyards[1858]}), .right({trees[1860], lumberyards[1860]}), .bottom_left({trees[1908], lumberyards[1908]}), .bottom({trees[1909], lumberyards[1909]}), .bottom_right({trees[1910], lumberyards[1910]}), .init(2'b00), .state({trees[1859], lumberyards[1859]}));
acre acre_37_10 (.clk(clk), .en(en), .top_left({trees[1809], lumberyards[1809]}), .top({trees[1810], lumberyards[1810]}), .top_right({trees[1811], lumberyards[1811]}), .left({trees[1859], lumberyards[1859]}), .right({trees[1861], lumberyards[1861]}), .bottom_left({trees[1909], lumberyards[1909]}), .bottom({trees[1910], lumberyards[1910]}), .bottom_right({trees[1911], lumberyards[1911]}), .init(2'b01), .state({trees[1860], lumberyards[1860]}));
acre acre_37_11 (.clk(clk), .en(en), .top_left({trees[1810], lumberyards[1810]}), .top({trees[1811], lumberyards[1811]}), .top_right({trees[1812], lumberyards[1812]}), .left({trees[1860], lumberyards[1860]}), .right({trees[1862], lumberyards[1862]}), .bottom_left({trees[1910], lumberyards[1910]}), .bottom({trees[1911], lumberyards[1911]}), .bottom_right({trees[1912], lumberyards[1912]}), .init(2'b10), .state({trees[1861], lumberyards[1861]}));
acre acre_37_12 (.clk(clk), .en(en), .top_left({trees[1811], lumberyards[1811]}), .top({trees[1812], lumberyards[1812]}), .top_right({trees[1813], lumberyards[1813]}), .left({trees[1861], lumberyards[1861]}), .right({trees[1863], lumberyards[1863]}), .bottom_left({trees[1911], lumberyards[1911]}), .bottom({trees[1912], lumberyards[1912]}), .bottom_right({trees[1913], lumberyards[1913]}), .init(2'b01), .state({trees[1862], lumberyards[1862]}));
acre acre_37_13 (.clk(clk), .en(en), .top_left({trees[1812], lumberyards[1812]}), .top({trees[1813], lumberyards[1813]}), .top_right({trees[1814], lumberyards[1814]}), .left({trees[1862], lumberyards[1862]}), .right({trees[1864], lumberyards[1864]}), .bottom_left({trees[1912], lumberyards[1912]}), .bottom({trees[1913], lumberyards[1913]}), .bottom_right({trees[1914], lumberyards[1914]}), .init(2'b01), .state({trees[1863], lumberyards[1863]}));
acre acre_37_14 (.clk(clk), .en(en), .top_left({trees[1813], lumberyards[1813]}), .top({trees[1814], lumberyards[1814]}), .top_right({trees[1815], lumberyards[1815]}), .left({trees[1863], lumberyards[1863]}), .right({trees[1865], lumberyards[1865]}), .bottom_left({trees[1913], lumberyards[1913]}), .bottom({trees[1914], lumberyards[1914]}), .bottom_right({trees[1915], lumberyards[1915]}), .init(2'b01), .state({trees[1864], lumberyards[1864]}));
acre acre_37_15 (.clk(clk), .en(en), .top_left({trees[1814], lumberyards[1814]}), .top({trees[1815], lumberyards[1815]}), .top_right({trees[1816], lumberyards[1816]}), .left({trees[1864], lumberyards[1864]}), .right({trees[1866], lumberyards[1866]}), .bottom_left({trees[1914], lumberyards[1914]}), .bottom({trees[1915], lumberyards[1915]}), .bottom_right({trees[1916], lumberyards[1916]}), .init(2'b10), .state({trees[1865], lumberyards[1865]}));
acre acre_37_16 (.clk(clk), .en(en), .top_left({trees[1815], lumberyards[1815]}), .top({trees[1816], lumberyards[1816]}), .top_right({trees[1817], lumberyards[1817]}), .left({trees[1865], lumberyards[1865]}), .right({trees[1867], lumberyards[1867]}), .bottom_left({trees[1915], lumberyards[1915]}), .bottom({trees[1916], lumberyards[1916]}), .bottom_right({trees[1917], lumberyards[1917]}), .init(2'b10), .state({trees[1866], lumberyards[1866]}));
acre acre_37_17 (.clk(clk), .en(en), .top_left({trees[1816], lumberyards[1816]}), .top({trees[1817], lumberyards[1817]}), .top_right({trees[1818], lumberyards[1818]}), .left({trees[1866], lumberyards[1866]}), .right({trees[1868], lumberyards[1868]}), .bottom_left({trees[1916], lumberyards[1916]}), .bottom({trees[1917], lumberyards[1917]}), .bottom_right({trees[1918], lumberyards[1918]}), .init(2'b00), .state({trees[1867], lumberyards[1867]}));
acre acre_37_18 (.clk(clk), .en(en), .top_left({trees[1817], lumberyards[1817]}), .top({trees[1818], lumberyards[1818]}), .top_right({trees[1819], lumberyards[1819]}), .left({trees[1867], lumberyards[1867]}), .right({trees[1869], lumberyards[1869]}), .bottom_left({trees[1917], lumberyards[1917]}), .bottom({trees[1918], lumberyards[1918]}), .bottom_right({trees[1919], lumberyards[1919]}), .init(2'b10), .state({trees[1868], lumberyards[1868]}));
acre acre_37_19 (.clk(clk), .en(en), .top_left({trees[1818], lumberyards[1818]}), .top({trees[1819], lumberyards[1819]}), .top_right({trees[1820], lumberyards[1820]}), .left({trees[1868], lumberyards[1868]}), .right({trees[1870], lumberyards[1870]}), .bottom_left({trees[1918], lumberyards[1918]}), .bottom({trees[1919], lumberyards[1919]}), .bottom_right({trees[1920], lumberyards[1920]}), .init(2'b10), .state({trees[1869], lumberyards[1869]}));
acre acre_37_20 (.clk(clk), .en(en), .top_left({trees[1819], lumberyards[1819]}), .top({trees[1820], lumberyards[1820]}), .top_right({trees[1821], lumberyards[1821]}), .left({trees[1869], lumberyards[1869]}), .right({trees[1871], lumberyards[1871]}), .bottom_left({trees[1919], lumberyards[1919]}), .bottom({trees[1920], lumberyards[1920]}), .bottom_right({trees[1921], lumberyards[1921]}), .init(2'b01), .state({trees[1870], lumberyards[1870]}));
acre acre_37_21 (.clk(clk), .en(en), .top_left({trees[1820], lumberyards[1820]}), .top({trees[1821], lumberyards[1821]}), .top_right({trees[1822], lumberyards[1822]}), .left({trees[1870], lumberyards[1870]}), .right({trees[1872], lumberyards[1872]}), .bottom_left({trees[1920], lumberyards[1920]}), .bottom({trees[1921], lumberyards[1921]}), .bottom_right({trees[1922], lumberyards[1922]}), .init(2'b01), .state({trees[1871], lumberyards[1871]}));
acre acre_37_22 (.clk(clk), .en(en), .top_left({trees[1821], lumberyards[1821]}), .top({trees[1822], lumberyards[1822]}), .top_right({trees[1823], lumberyards[1823]}), .left({trees[1871], lumberyards[1871]}), .right({trees[1873], lumberyards[1873]}), .bottom_left({trees[1921], lumberyards[1921]}), .bottom({trees[1922], lumberyards[1922]}), .bottom_right({trees[1923], lumberyards[1923]}), .init(2'b01), .state({trees[1872], lumberyards[1872]}));
acre acre_37_23 (.clk(clk), .en(en), .top_left({trees[1822], lumberyards[1822]}), .top({trees[1823], lumberyards[1823]}), .top_right({trees[1824], lumberyards[1824]}), .left({trees[1872], lumberyards[1872]}), .right({trees[1874], lumberyards[1874]}), .bottom_left({trees[1922], lumberyards[1922]}), .bottom({trees[1923], lumberyards[1923]}), .bottom_right({trees[1924], lumberyards[1924]}), .init(2'b10), .state({trees[1873], lumberyards[1873]}));
acre acre_37_24 (.clk(clk), .en(en), .top_left({trees[1823], lumberyards[1823]}), .top({trees[1824], lumberyards[1824]}), .top_right({trees[1825], lumberyards[1825]}), .left({trees[1873], lumberyards[1873]}), .right({trees[1875], lumberyards[1875]}), .bottom_left({trees[1923], lumberyards[1923]}), .bottom({trees[1924], lumberyards[1924]}), .bottom_right({trees[1925], lumberyards[1925]}), .init(2'b00), .state({trees[1874], lumberyards[1874]}));
acre acre_37_25 (.clk(clk), .en(en), .top_left({trees[1824], lumberyards[1824]}), .top({trees[1825], lumberyards[1825]}), .top_right({trees[1826], lumberyards[1826]}), .left({trees[1874], lumberyards[1874]}), .right({trees[1876], lumberyards[1876]}), .bottom_left({trees[1924], lumberyards[1924]}), .bottom({trees[1925], lumberyards[1925]}), .bottom_right({trees[1926], lumberyards[1926]}), .init(2'b00), .state({trees[1875], lumberyards[1875]}));
acre acre_37_26 (.clk(clk), .en(en), .top_left({trees[1825], lumberyards[1825]}), .top({trees[1826], lumberyards[1826]}), .top_right({trees[1827], lumberyards[1827]}), .left({trees[1875], lumberyards[1875]}), .right({trees[1877], lumberyards[1877]}), .bottom_left({trees[1925], lumberyards[1925]}), .bottom({trees[1926], lumberyards[1926]}), .bottom_right({trees[1927], lumberyards[1927]}), .init(2'b10), .state({trees[1876], lumberyards[1876]}));
acre acre_37_27 (.clk(clk), .en(en), .top_left({trees[1826], lumberyards[1826]}), .top({trees[1827], lumberyards[1827]}), .top_right({trees[1828], lumberyards[1828]}), .left({trees[1876], lumberyards[1876]}), .right({trees[1878], lumberyards[1878]}), .bottom_left({trees[1926], lumberyards[1926]}), .bottom({trees[1927], lumberyards[1927]}), .bottom_right({trees[1928], lumberyards[1928]}), .init(2'b00), .state({trees[1877], lumberyards[1877]}));
acre acre_37_28 (.clk(clk), .en(en), .top_left({trees[1827], lumberyards[1827]}), .top({trees[1828], lumberyards[1828]}), .top_right({trees[1829], lumberyards[1829]}), .left({trees[1877], lumberyards[1877]}), .right({trees[1879], lumberyards[1879]}), .bottom_left({trees[1927], lumberyards[1927]}), .bottom({trees[1928], lumberyards[1928]}), .bottom_right({trees[1929], lumberyards[1929]}), .init(2'b00), .state({trees[1878], lumberyards[1878]}));
acre acre_37_29 (.clk(clk), .en(en), .top_left({trees[1828], lumberyards[1828]}), .top({trees[1829], lumberyards[1829]}), .top_right({trees[1830], lumberyards[1830]}), .left({trees[1878], lumberyards[1878]}), .right({trees[1880], lumberyards[1880]}), .bottom_left({trees[1928], lumberyards[1928]}), .bottom({trees[1929], lumberyards[1929]}), .bottom_right({trees[1930], lumberyards[1930]}), .init(2'b01), .state({trees[1879], lumberyards[1879]}));
acre acre_37_30 (.clk(clk), .en(en), .top_left({trees[1829], lumberyards[1829]}), .top({trees[1830], lumberyards[1830]}), .top_right({trees[1831], lumberyards[1831]}), .left({trees[1879], lumberyards[1879]}), .right({trees[1881], lumberyards[1881]}), .bottom_left({trees[1929], lumberyards[1929]}), .bottom({trees[1930], lumberyards[1930]}), .bottom_right({trees[1931], lumberyards[1931]}), .init(2'b00), .state({trees[1880], lumberyards[1880]}));
acre acre_37_31 (.clk(clk), .en(en), .top_left({trees[1830], lumberyards[1830]}), .top({trees[1831], lumberyards[1831]}), .top_right({trees[1832], lumberyards[1832]}), .left({trees[1880], lumberyards[1880]}), .right({trees[1882], lumberyards[1882]}), .bottom_left({trees[1930], lumberyards[1930]}), .bottom({trees[1931], lumberyards[1931]}), .bottom_right({trees[1932], lumberyards[1932]}), .init(2'b10), .state({trees[1881], lumberyards[1881]}));
acre acre_37_32 (.clk(clk), .en(en), .top_left({trees[1831], lumberyards[1831]}), .top({trees[1832], lumberyards[1832]}), .top_right({trees[1833], lumberyards[1833]}), .left({trees[1881], lumberyards[1881]}), .right({trees[1883], lumberyards[1883]}), .bottom_left({trees[1931], lumberyards[1931]}), .bottom({trees[1932], lumberyards[1932]}), .bottom_right({trees[1933], lumberyards[1933]}), .init(2'b01), .state({trees[1882], lumberyards[1882]}));
acre acre_37_33 (.clk(clk), .en(en), .top_left({trees[1832], lumberyards[1832]}), .top({trees[1833], lumberyards[1833]}), .top_right({trees[1834], lumberyards[1834]}), .left({trees[1882], lumberyards[1882]}), .right({trees[1884], lumberyards[1884]}), .bottom_left({trees[1932], lumberyards[1932]}), .bottom({trees[1933], lumberyards[1933]}), .bottom_right({trees[1934], lumberyards[1934]}), .init(2'b00), .state({trees[1883], lumberyards[1883]}));
acre acre_37_34 (.clk(clk), .en(en), .top_left({trees[1833], lumberyards[1833]}), .top({trees[1834], lumberyards[1834]}), .top_right({trees[1835], lumberyards[1835]}), .left({trees[1883], lumberyards[1883]}), .right({trees[1885], lumberyards[1885]}), .bottom_left({trees[1933], lumberyards[1933]}), .bottom({trees[1934], lumberyards[1934]}), .bottom_right({trees[1935], lumberyards[1935]}), .init(2'b00), .state({trees[1884], lumberyards[1884]}));
acre acre_37_35 (.clk(clk), .en(en), .top_left({trees[1834], lumberyards[1834]}), .top({trees[1835], lumberyards[1835]}), .top_right({trees[1836], lumberyards[1836]}), .left({trees[1884], lumberyards[1884]}), .right({trees[1886], lumberyards[1886]}), .bottom_left({trees[1934], lumberyards[1934]}), .bottom({trees[1935], lumberyards[1935]}), .bottom_right({trees[1936], lumberyards[1936]}), .init(2'b00), .state({trees[1885], lumberyards[1885]}));
acre acre_37_36 (.clk(clk), .en(en), .top_left({trees[1835], lumberyards[1835]}), .top({trees[1836], lumberyards[1836]}), .top_right({trees[1837], lumberyards[1837]}), .left({trees[1885], lumberyards[1885]}), .right({trees[1887], lumberyards[1887]}), .bottom_left({trees[1935], lumberyards[1935]}), .bottom({trees[1936], lumberyards[1936]}), .bottom_right({trees[1937], lumberyards[1937]}), .init(2'b00), .state({trees[1886], lumberyards[1886]}));
acre acre_37_37 (.clk(clk), .en(en), .top_left({trees[1836], lumberyards[1836]}), .top({trees[1837], lumberyards[1837]}), .top_right({trees[1838], lumberyards[1838]}), .left({trees[1886], lumberyards[1886]}), .right({trees[1888], lumberyards[1888]}), .bottom_left({trees[1936], lumberyards[1936]}), .bottom({trees[1937], lumberyards[1937]}), .bottom_right({trees[1938], lumberyards[1938]}), .init(2'b10), .state({trees[1887], lumberyards[1887]}));
acre acre_37_38 (.clk(clk), .en(en), .top_left({trees[1837], lumberyards[1837]}), .top({trees[1838], lumberyards[1838]}), .top_right({trees[1839], lumberyards[1839]}), .left({trees[1887], lumberyards[1887]}), .right({trees[1889], lumberyards[1889]}), .bottom_left({trees[1937], lumberyards[1937]}), .bottom({trees[1938], lumberyards[1938]}), .bottom_right({trees[1939], lumberyards[1939]}), .init(2'b01), .state({trees[1888], lumberyards[1888]}));
acre acre_37_39 (.clk(clk), .en(en), .top_left({trees[1838], lumberyards[1838]}), .top({trees[1839], lumberyards[1839]}), .top_right({trees[1840], lumberyards[1840]}), .left({trees[1888], lumberyards[1888]}), .right({trees[1890], lumberyards[1890]}), .bottom_left({trees[1938], lumberyards[1938]}), .bottom({trees[1939], lumberyards[1939]}), .bottom_right({trees[1940], lumberyards[1940]}), .init(2'b00), .state({trees[1889], lumberyards[1889]}));
acre acre_37_40 (.clk(clk), .en(en), .top_left({trees[1839], lumberyards[1839]}), .top({trees[1840], lumberyards[1840]}), .top_right({trees[1841], lumberyards[1841]}), .left({trees[1889], lumberyards[1889]}), .right({trees[1891], lumberyards[1891]}), .bottom_left({trees[1939], lumberyards[1939]}), .bottom({trees[1940], lumberyards[1940]}), .bottom_right({trees[1941], lumberyards[1941]}), .init(2'b00), .state({trees[1890], lumberyards[1890]}));
acre acre_37_41 (.clk(clk), .en(en), .top_left({trees[1840], lumberyards[1840]}), .top({trees[1841], lumberyards[1841]}), .top_right({trees[1842], lumberyards[1842]}), .left({trees[1890], lumberyards[1890]}), .right({trees[1892], lumberyards[1892]}), .bottom_left({trees[1940], lumberyards[1940]}), .bottom({trees[1941], lumberyards[1941]}), .bottom_right({trees[1942], lumberyards[1942]}), .init(2'b00), .state({trees[1891], lumberyards[1891]}));
acre acre_37_42 (.clk(clk), .en(en), .top_left({trees[1841], lumberyards[1841]}), .top({trees[1842], lumberyards[1842]}), .top_right({trees[1843], lumberyards[1843]}), .left({trees[1891], lumberyards[1891]}), .right({trees[1893], lumberyards[1893]}), .bottom_left({trees[1941], lumberyards[1941]}), .bottom({trees[1942], lumberyards[1942]}), .bottom_right({trees[1943], lumberyards[1943]}), .init(2'b00), .state({trees[1892], lumberyards[1892]}));
acre acre_37_43 (.clk(clk), .en(en), .top_left({trees[1842], lumberyards[1842]}), .top({trees[1843], lumberyards[1843]}), .top_right({trees[1844], lumberyards[1844]}), .left({trees[1892], lumberyards[1892]}), .right({trees[1894], lumberyards[1894]}), .bottom_left({trees[1942], lumberyards[1942]}), .bottom({trees[1943], lumberyards[1943]}), .bottom_right({trees[1944], lumberyards[1944]}), .init(2'b10), .state({trees[1893], lumberyards[1893]}));
acre acre_37_44 (.clk(clk), .en(en), .top_left({trees[1843], lumberyards[1843]}), .top({trees[1844], lumberyards[1844]}), .top_right({trees[1845], lumberyards[1845]}), .left({trees[1893], lumberyards[1893]}), .right({trees[1895], lumberyards[1895]}), .bottom_left({trees[1943], lumberyards[1943]}), .bottom({trees[1944], lumberyards[1944]}), .bottom_right({trees[1945], lumberyards[1945]}), .init(2'b00), .state({trees[1894], lumberyards[1894]}));
acre acre_37_45 (.clk(clk), .en(en), .top_left({trees[1844], lumberyards[1844]}), .top({trees[1845], lumberyards[1845]}), .top_right({trees[1846], lumberyards[1846]}), .left({trees[1894], lumberyards[1894]}), .right({trees[1896], lumberyards[1896]}), .bottom_left({trees[1944], lumberyards[1944]}), .bottom({trees[1945], lumberyards[1945]}), .bottom_right({trees[1946], lumberyards[1946]}), .init(2'b01), .state({trees[1895], lumberyards[1895]}));
acre acre_37_46 (.clk(clk), .en(en), .top_left({trees[1845], lumberyards[1845]}), .top({trees[1846], lumberyards[1846]}), .top_right({trees[1847], lumberyards[1847]}), .left({trees[1895], lumberyards[1895]}), .right({trees[1897], lumberyards[1897]}), .bottom_left({trees[1945], lumberyards[1945]}), .bottom({trees[1946], lumberyards[1946]}), .bottom_right({trees[1947], lumberyards[1947]}), .init(2'b00), .state({trees[1896], lumberyards[1896]}));
acre acre_37_47 (.clk(clk), .en(en), .top_left({trees[1846], lumberyards[1846]}), .top({trees[1847], lumberyards[1847]}), .top_right({trees[1848], lumberyards[1848]}), .left({trees[1896], lumberyards[1896]}), .right({trees[1898], lumberyards[1898]}), .bottom_left({trees[1946], lumberyards[1946]}), .bottom({trees[1947], lumberyards[1947]}), .bottom_right({trees[1948], lumberyards[1948]}), .init(2'b10), .state({trees[1897], lumberyards[1897]}));
acre acre_37_48 (.clk(clk), .en(en), .top_left({trees[1847], lumberyards[1847]}), .top({trees[1848], lumberyards[1848]}), .top_right({trees[1849], lumberyards[1849]}), .left({trees[1897], lumberyards[1897]}), .right({trees[1899], lumberyards[1899]}), .bottom_left({trees[1947], lumberyards[1947]}), .bottom({trees[1948], lumberyards[1948]}), .bottom_right({trees[1949], lumberyards[1949]}), .init(2'b00), .state({trees[1898], lumberyards[1898]}));
acre acre_37_49 (.clk(clk), .en(en), .top_left({trees[1848], lumberyards[1848]}), .top({trees[1849], lumberyards[1849]}), .top_right(2'b0), .left({trees[1898], lumberyards[1898]}), .right(2'b0), .bottom_left({trees[1948], lumberyards[1948]}), .bottom({trees[1949], lumberyards[1949]}), .bottom_right(2'b0), .init(2'b00), .state({trees[1899], lumberyards[1899]}));
acre acre_38_0 (.clk(clk), .en(en), .top_left(2'b0), .top({trees[1850], lumberyards[1850]}), .top_right({trees[1851], lumberyards[1851]}), .left(2'b0), .right({trees[1901], lumberyards[1901]}), .bottom_left(2'b0), .bottom({trees[1950], lumberyards[1950]}), .bottom_right({trees[1951], lumberyards[1951]}), .init(2'b00), .state({trees[1900], lumberyards[1900]}));
acre acre_38_1 (.clk(clk), .en(en), .top_left({trees[1850], lumberyards[1850]}), .top({trees[1851], lumberyards[1851]}), .top_right({trees[1852], lumberyards[1852]}), .left({trees[1900], lumberyards[1900]}), .right({trees[1902], lumberyards[1902]}), .bottom_left({trees[1950], lumberyards[1950]}), .bottom({trees[1951], lumberyards[1951]}), .bottom_right({trees[1952], lumberyards[1952]}), .init(2'b10), .state({trees[1901], lumberyards[1901]}));
acre acre_38_2 (.clk(clk), .en(en), .top_left({trees[1851], lumberyards[1851]}), .top({trees[1852], lumberyards[1852]}), .top_right({trees[1853], lumberyards[1853]}), .left({trees[1901], lumberyards[1901]}), .right({trees[1903], lumberyards[1903]}), .bottom_left({trees[1951], lumberyards[1951]}), .bottom({trees[1952], lumberyards[1952]}), .bottom_right({trees[1953], lumberyards[1953]}), .init(2'b10), .state({trees[1902], lumberyards[1902]}));
acre acre_38_3 (.clk(clk), .en(en), .top_left({trees[1852], lumberyards[1852]}), .top({trees[1853], lumberyards[1853]}), .top_right({trees[1854], lumberyards[1854]}), .left({trees[1902], lumberyards[1902]}), .right({trees[1904], lumberyards[1904]}), .bottom_left({trees[1952], lumberyards[1952]}), .bottom({trees[1953], lumberyards[1953]}), .bottom_right({trees[1954], lumberyards[1954]}), .init(2'b00), .state({trees[1903], lumberyards[1903]}));
acre acre_38_4 (.clk(clk), .en(en), .top_left({trees[1853], lumberyards[1853]}), .top({trees[1854], lumberyards[1854]}), .top_right({trees[1855], lumberyards[1855]}), .left({trees[1903], lumberyards[1903]}), .right({trees[1905], lumberyards[1905]}), .bottom_left({trees[1953], lumberyards[1953]}), .bottom({trees[1954], lumberyards[1954]}), .bottom_right({trees[1955], lumberyards[1955]}), .init(2'b00), .state({trees[1904], lumberyards[1904]}));
acre acre_38_5 (.clk(clk), .en(en), .top_left({trees[1854], lumberyards[1854]}), .top({trees[1855], lumberyards[1855]}), .top_right({trees[1856], lumberyards[1856]}), .left({trees[1904], lumberyards[1904]}), .right({trees[1906], lumberyards[1906]}), .bottom_left({trees[1954], lumberyards[1954]}), .bottom({trees[1955], lumberyards[1955]}), .bottom_right({trees[1956], lumberyards[1956]}), .init(2'b10), .state({trees[1905], lumberyards[1905]}));
acre acre_38_6 (.clk(clk), .en(en), .top_left({trees[1855], lumberyards[1855]}), .top({trees[1856], lumberyards[1856]}), .top_right({trees[1857], lumberyards[1857]}), .left({trees[1905], lumberyards[1905]}), .right({trees[1907], lumberyards[1907]}), .bottom_left({trees[1955], lumberyards[1955]}), .bottom({trees[1956], lumberyards[1956]}), .bottom_right({trees[1957], lumberyards[1957]}), .init(2'b01), .state({trees[1906], lumberyards[1906]}));
acre acre_38_7 (.clk(clk), .en(en), .top_left({trees[1856], lumberyards[1856]}), .top({trees[1857], lumberyards[1857]}), .top_right({trees[1858], lumberyards[1858]}), .left({trees[1906], lumberyards[1906]}), .right({trees[1908], lumberyards[1908]}), .bottom_left({trees[1956], lumberyards[1956]}), .bottom({trees[1957], lumberyards[1957]}), .bottom_right({trees[1958], lumberyards[1958]}), .init(2'b00), .state({trees[1907], lumberyards[1907]}));
acre acre_38_8 (.clk(clk), .en(en), .top_left({trees[1857], lumberyards[1857]}), .top({trees[1858], lumberyards[1858]}), .top_right({trees[1859], lumberyards[1859]}), .left({trees[1907], lumberyards[1907]}), .right({trees[1909], lumberyards[1909]}), .bottom_left({trees[1957], lumberyards[1957]}), .bottom({trees[1958], lumberyards[1958]}), .bottom_right({trees[1959], lumberyards[1959]}), .init(2'b00), .state({trees[1908], lumberyards[1908]}));
acre acre_38_9 (.clk(clk), .en(en), .top_left({trees[1858], lumberyards[1858]}), .top({trees[1859], lumberyards[1859]}), .top_right({trees[1860], lumberyards[1860]}), .left({trees[1908], lumberyards[1908]}), .right({trees[1910], lumberyards[1910]}), .bottom_left({trees[1958], lumberyards[1958]}), .bottom({trees[1959], lumberyards[1959]}), .bottom_right({trees[1960], lumberyards[1960]}), .init(2'b00), .state({trees[1909], lumberyards[1909]}));
acre acre_38_10 (.clk(clk), .en(en), .top_left({trees[1859], lumberyards[1859]}), .top({trees[1860], lumberyards[1860]}), .top_right({trees[1861], lumberyards[1861]}), .left({trees[1909], lumberyards[1909]}), .right({trees[1911], lumberyards[1911]}), .bottom_left({trees[1959], lumberyards[1959]}), .bottom({trees[1960], lumberyards[1960]}), .bottom_right({trees[1961], lumberyards[1961]}), .init(2'b00), .state({trees[1910], lumberyards[1910]}));
acre acre_38_11 (.clk(clk), .en(en), .top_left({trees[1860], lumberyards[1860]}), .top({trees[1861], lumberyards[1861]}), .top_right({trees[1862], lumberyards[1862]}), .left({trees[1910], lumberyards[1910]}), .right({trees[1912], lumberyards[1912]}), .bottom_left({trees[1960], lumberyards[1960]}), .bottom({trees[1961], lumberyards[1961]}), .bottom_right({trees[1962], lumberyards[1962]}), .init(2'b01), .state({trees[1911], lumberyards[1911]}));
acre acre_38_12 (.clk(clk), .en(en), .top_left({trees[1861], lumberyards[1861]}), .top({trees[1862], lumberyards[1862]}), .top_right({trees[1863], lumberyards[1863]}), .left({trees[1911], lumberyards[1911]}), .right({trees[1913], lumberyards[1913]}), .bottom_left({trees[1961], lumberyards[1961]}), .bottom({trees[1962], lumberyards[1962]}), .bottom_right({trees[1963], lumberyards[1963]}), .init(2'b01), .state({trees[1912], lumberyards[1912]}));
acre acre_38_13 (.clk(clk), .en(en), .top_left({trees[1862], lumberyards[1862]}), .top({trees[1863], lumberyards[1863]}), .top_right({trees[1864], lumberyards[1864]}), .left({trees[1912], lumberyards[1912]}), .right({trees[1914], lumberyards[1914]}), .bottom_left({trees[1962], lumberyards[1962]}), .bottom({trees[1963], lumberyards[1963]}), .bottom_right({trees[1964], lumberyards[1964]}), .init(2'b01), .state({trees[1913], lumberyards[1913]}));
acre acre_38_14 (.clk(clk), .en(en), .top_left({trees[1863], lumberyards[1863]}), .top({trees[1864], lumberyards[1864]}), .top_right({trees[1865], lumberyards[1865]}), .left({trees[1913], lumberyards[1913]}), .right({trees[1915], lumberyards[1915]}), .bottom_left({trees[1963], lumberyards[1963]}), .bottom({trees[1964], lumberyards[1964]}), .bottom_right({trees[1965], lumberyards[1965]}), .init(2'b00), .state({trees[1914], lumberyards[1914]}));
acre acre_38_15 (.clk(clk), .en(en), .top_left({trees[1864], lumberyards[1864]}), .top({trees[1865], lumberyards[1865]}), .top_right({trees[1866], lumberyards[1866]}), .left({trees[1914], lumberyards[1914]}), .right({trees[1916], lumberyards[1916]}), .bottom_left({trees[1964], lumberyards[1964]}), .bottom({trees[1965], lumberyards[1965]}), .bottom_right({trees[1966], lumberyards[1966]}), .init(2'b10), .state({trees[1915], lumberyards[1915]}));
acre acre_38_16 (.clk(clk), .en(en), .top_left({trees[1865], lumberyards[1865]}), .top({trees[1866], lumberyards[1866]}), .top_right({trees[1867], lumberyards[1867]}), .left({trees[1915], lumberyards[1915]}), .right({trees[1917], lumberyards[1917]}), .bottom_left({trees[1965], lumberyards[1965]}), .bottom({trees[1966], lumberyards[1966]}), .bottom_right({trees[1967], lumberyards[1967]}), .init(2'b10), .state({trees[1916], lumberyards[1916]}));
acre acre_38_17 (.clk(clk), .en(en), .top_left({trees[1866], lumberyards[1866]}), .top({trees[1867], lumberyards[1867]}), .top_right({trees[1868], lumberyards[1868]}), .left({trees[1916], lumberyards[1916]}), .right({trees[1918], lumberyards[1918]}), .bottom_left({trees[1966], lumberyards[1966]}), .bottom({trees[1967], lumberyards[1967]}), .bottom_right({trees[1968], lumberyards[1968]}), .init(2'b01), .state({trees[1917], lumberyards[1917]}));
acre acre_38_18 (.clk(clk), .en(en), .top_left({trees[1867], lumberyards[1867]}), .top({trees[1868], lumberyards[1868]}), .top_right({trees[1869], lumberyards[1869]}), .left({trees[1917], lumberyards[1917]}), .right({trees[1919], lumberyards[1919]}), .bottom_left({trees[1967], lumberyards[1967]}), .bottom({trees[1968], lumberyards[1968]}), .bottom_right({trees[1969], lumberyards[1969]}), .init(2'b00), .state({trees[1918], lumberyards[1918]}));
acre acre_38_19 (.clk(clk), .en(en), .top_left({trees[1868], lumberyards[1868]}), .top({trees[1869], lumberyards[1869]}), .top_right({trees[1870], lumberyards[1870]}), .left({trees[1918], lumberyards[1918]}), .right({trees[1920], lumberyards[1920]}), .bottom_left({trees[1968], lumberyards[1968]}), .bottom({trees[1969], lumberyards[1969]}), .bottom_right({trees[1970], lumberyards[1970]}), .init(2'b00), .state({trees[1919], lumberyards[1919]}));
acre acre_38_20 (.clk(clk), .en(en), .top_left({trees[1869], lumberyards[1869]}), .top({trees[1870], lumberyards[1870]}), .top_right({trees[1871], lumberyards[1871]}), .left({trees[1919], lumberyards[1919]}), .right({trees[1921], lumberyards[1921]}), .bottom_left({trees[1969], lumberyards[1969]}), .bottom({trees[1970], lumberyards[1970]}), .bottom_right({trees[1971], lumberyards[1971]}), .init(2'b01), .state({trees[1920], lumberyards[1920]}));
acre acre_38_21 (.clk(clk), .en(en), .top_left({trees[1870], lumberyards[1870]}), .top({trees[1871], lumberyards[1871]}), .top_right({trees[1872], lumberyards[1872]}), .left({trees[1920], lumberyards[1920]}), .right({trees[1922], lumberyards[1922]}), .bottom_left({trees[1970], lumberyards[1970]}), .bottom({trees[1971], lumberyards[1971]}), .bottom_right({trees[1972], lumberyards[1972]}), .init(2'b00), .state({trees[1921], lumberyards[1921]}));
acre acre_38_22 (.clk(clk), .en(en), .top_left({trees[1871], lumberyards[1871]}), .top({trees[1872], lumberyards[1872]}), .top_right({trees[1873], lumberyards[1873]}), .left({trees[1921], lumberyards[1921]}), .right({trees[1923], lumberyards[1923]}), .bottom_left({trees[1971], lumberyards[1971]}), .bottom({trees[1972], lumberyards[1972]}), .bottom_right({trees[1973], lumberyards[1973]}), .init(2'b10), .state({trees[1922], lumberyards[1922]}));
acre acre_38_23 (.clk(clk), .en(en), .top_left({trees[1872], lumberyards[1872]}), .top({trees[1873], lumberyards[1873]}), .top_right({trees[1874], lumberyards[1874]}), .left({trees[1922], lumberyards[1922]}), .right({trees[1924], lumberyards[1924]}), .bottom_left({trees[1972], lumberyards[1972]}), .bottom({trees[1973], lumberyards[1973]}), .bottom_right({trees[1974], lumberyards[1974]}), .init(2'b00), .state({trees[1923], lumberyards[1923]}));
acre acre_38_24 (.clk(clk), .en(en), .top_left({trees[1873], lumberyards[1873]}), .top({trees[1874], lumberyards[1874]}), .top_right({trees[1875], lumberyards[1875]}), .left({trees[1923], lumberyards[1923]}), .right({trees[1925], lumberyards[1925]}), .bottom_left({trees[1973], lumberyards[1973]}), .bottom({trees[1974], lumberyards[1974]}), .bottom_right({trees[1975], lumberyards[1975]}), .init(2'b00), .state({trees[1924], lumberyards[1924]}));
acre acre_38_25 (.clk(clk), .en(en), .top_left({trees[1874], lumberyards[1874]}), .top({trees[1875], lumberyards[1875]}), .top_right({trees[1876], lumberyards[1876]}), .left({trees[1924], lumberyards[1924]}), .right({trees[1926], lumberyards[1926]}), .bottom_left({trees[1974], lumberyards[1974]}), .bottom({trees[1975], lumberyards[1975]}), .bottom_right({trees[1976], lumberyards[1976]}), .init(2'b00), .state({trees[1925], lumberyards[1925]}));
acre acre_38_26 (.clk(clk), .en(en), .top_left({trees[1875], lumberyards[1875]}), .top({trees[1876], lumberyards[1876]}), .top_right({trees[1877], lumberyards[1877]}), .left({trees[1925], lumberyards[1925]}), .right({trees[1927], lumberyards[1927]}), .bottom_left({trees[1975], lumberyards[1975]}), .bottom({trees[1976], lumberyards[1976]}), .bottom_right({trees[1977], lumberyards[1977]}), .init(2'b00), .state({trees[1926], lumberyards[1926]}));
acre acre_38_27 (.clk(clk), .en(en), .top_left({trees[1876], lumberyards[1876]}), .top({trees[1877], lumberyards[1877]}), .top_right({trees[1878], lumberyards[1878]}), .left({trees[1926], lumberyards[1926]}), .right({trees[1928], lumberyards[1928]}), .bottom_left({trees[1976], lumberyards[1976]}), .bottom({trees[1977], lumberyards[1977]}), .bottom_right({trees[1978], lumberyards[1978]}), .init(2'b00), .state({trees[1927], lumberyards[1927]}));
acre acre_38_28 (.clk(clk), .en(en), .top_left({trees[1877], lumberyards[1877]}), .top({trees[1878], lumberyards[1878]}), .top_right({trees[1879], lumberyards[1879]}), .left({trees[1927], lumberyards[1927]}), .right({trees[1929], lumberyards[1929]}), .bottom_left({trees[1977], lumberyards[1977]}), .bottom({trees[1978], lumberyards[1978]}), .bottom_right({trees[1979], lumberyards[1979]}), .init(2'b00), .state({trees[1928], lumberyards[1928]}));
acre acre_38_29 (.clk(clk), .en(en), .top_left({trees[1878], lumberyards[1878]}), .top({trees[1879], lumberyards[1879]}), .top_right({trees[1880], lumberyards[1880]}), .left({trees[1928], lumberyards[1928]}), .right({trees[1930], lumberyards[1930]}), .bottom_left({trees[1978], lumberyards[1978]}), .bottom({trees[1979], lumberyards[1979]}), .bottom_right({trees[1980], lumberyards[1980]}), .init(2'b00), .state({trees[1929], lumberyards[1929]}));
acre acre_38_30 (.clk(clk), .en(en), .top_left({trees[1879], lumberyards[1879]}), .top({trees[1880], lumberyards[1880]}), .top_right({trees[1881], lumberyards[1881]}), .left({trees[1929], lumberyards[1929]}), .right({trees[1931], lumberyards[1931]}), .bottom_left({trees[1979], lumberyards[1979]}), .bottom({trees[1980], lumberyards[1980]}), .bottom_right({trees[1981], lumberyards[1981]}), .init(2'b00), .state({trees[1930], lumberyards[1930]}));
acre acre_38_31 (.clk(clk), .en(en), .top_left({trees[1880], lumberyards[1880]}), .top({trees[1881], lumberyards[1881]}), .top_right({trees[1882], lumberyards[1882]}), .left({trees[1930], lumberyards[1930]}), .right({trees[1932], lumberyards[1932]}), .bottom_left({trees[1980], lumberyards[1980]}), .bottom({trees[1981], lumberyards[1981]}), .bottom_right({trees[1982], lumberyards[1982]}), .init(2'b01), .state({trees[1931], lumberyards[1931]}));
acre acre_38_32 (.clk(clk), .en(en), .top_left({trees[1881], lumberyards[1881]}), .top({trees[1882], lumberyards[1882]}), .top_right({trees[1883], lumberyards[1883]}), .left({trees[1931], lumberyards[1931]}), .right({trees[1933], lumberyards[1933]}), .bottom_left({trees[1981], lumberyards[1981]}), .bottom({trees[1982], lumberyards[1982]}), .bottom_right({trees[1983], lumberyards[1983]}), .init(2'b01), .state({trees[1932], lumberyards[1932]}));
acre acre_38_33 (.clk(clk), .en(en), .top_left({trees[1882], lumberyards[1882]}), .top({trees[1883], lumberyards[1883]}), .top_right({trees[1884], lumberyards[1884]}), .left({trees[1932], lumberyards[1932]}), .right({trees[1934], lumberyards[1934]}), .bottom_left({trees[1982], lumberyards[1982]}), .bottom({trees[1983], lumberyards[1983]}), .bottom_right({trees[1984], lumberyards[1984]}), .init(2'b01), .state({trees[1933], lumberyards[1933]}));
acre acre_38_34 (.clk(clk), .en(en), .top_left({trees[1883], lumberyards[1883]}), .top({trees[1884], lumberyards[1884]}), .top_right({trees[1885], lumberyards[1885]}), .left({trees[1933], lumberyards[1933]}), .right({trees[1935], lumberyards[1935]}), .bottom_left({trees[1983], lumberyards[1983]}), .bottom({trees[1984], lumberyards[1984]}), .bottom_right({trees[1985], lumberyards[1985]}), .init(2'b00), .state({trees[1934], lumberyards[1934]}));
acre acre_38_35 (.clk(clk), .en(en), .top_left({trees[1884], lumberyards[1884]}), .top({trees[1885], lumberyards[1885]}), .top_right({trees[1886], lumberyards[1886]}), .left({trees[1934], lumberyards[1934]}), .right({trees[1936], lumberyards[1936]}), .bottom_left({trees[1984], lumberyards[1984]}), .bottom({trees[1985], lumberyards[1985]}), .bottom_right({trees[1986], lumberyards[1986]}), .init(2'b00), .state({trees[1935], lumberyards[1935]}));
acre acre_38_36 (.clk(clk), .en(en), .top_left({trees[1885], lumberyards[1885]}), .top({trees[1886], lumberyards[1886]}), .top_right({trees[1887], lumberyards[1887]}), .left({trees[1935], lumberyards[1935]}), .right({trees[1937], lumberyards[1937]}), .bottom_left({trees[1985], lumberyards[1985]}), .bottom({trees[1986], lumberyards[1986]}), .bottom_right({trees[1987], lumberyards[1987]}), .init(2'b10), .state({trees[1936], lumberyards[1936]}));
acre acre_38_37 (.clk(clk), .en(en), .top_left({trees[1886], lumberyards[1886]}), .top({trees[1887], lumberyards[1887]}), .top_right({trees[1888], lumberyards[1888]}), .left({trees[1936], lumberyards[1936]}), .right({trees[1938], lumberyards[1938]}), .bottom_left({trees[1986], lumberyards[1986]}), .bottom({trees[1987], lumberyards[1987]}), .bottom_right({trees[1988], lumberyards[1988]}), .init(2'b00), .state({trees[1937], lumberyards[1937]}));
acre acre_38_38 (.clk(clk), .en(en), .top_left({trees[1887], lumberyards[1887]}), .top({trees[1888], lumberyards[1888]}), .top_right({trees[1889], lumberyards[1889]}), .left({trees[1937], lumberyards[1937]}), .right({trees[1939], lumberyards[1939]}), .bottom_left({trees[1987], lumberyards[1987]}), .bottom({trees[1988], lumberyards[1988]}), .bottom_right({trees[1989], lumberyards[1989]}), .init(2'b01), .state({trees[1938], lumberyards[1938]}));
acre acre_38_39 (.clk(clk), .en(en), .top_left({trees[1888], lumberyards[1888]}), .top({trees[1889], lumberyards[1889]}), .top_right({trees[1890], lumberyards[1890]}), .left({trees[1938], lumberyards[1938]}), .right({trees[1940], lumberyards[1940]}), .bottom_left({trees[1988], lumberyards[1988]}), .bottom({trees[1989], lumberyards[1989]}), .bottom_right({trees[1990], lumberyards[1990]}), .init(2'b00), .state({trees[1939], lumberyards[1939]}));
acre acre_38_40 (.clk(clk), .en(en), .top_left({trees[1889], lumberyards[1889]}), .top({trees[1890], lumberyards[1890]}), .top_right({trees[1891], lumberyards[1891]}), .left({trees[1939], lumberyards[1939]}), .right({trees[1941], lumberyards[1941]}), .bottom_left({trees[1989], lumberyards[1989]}), .bottom({trees[1990], lumberyards[1990]}), .bottom_right({trees[1991], lumberyards[1991]}), .init(2'b00), .state({trees[1940], lumberyards[1940]}));
acre acre_38_41 (.clk(clk), .en(en), .top_left({trees[1890], lumberyards[1890]}), .top({trees[1891], lumberyards[1891]}), .top_right({trees[1892], lumberyards[1892]}), .left({trees[1940], lumberyards[1940]}), .right({trees[1942], lumberyards[1942]}), .bottom_left({trees[1990], lumberyards[1990]}), .bottom({trees[1991], lumberyards[1991]}), .bottom_right({trees[1992], lumberyards[1992]}), .init(2'b00), .state({trees[1941], lumberyards[1941]}));
acre acre_38_42 (.clk(clk), .en(en), .top_left({trees[1891], lumberyards[1891]}), .top({trees[1892], lumberyards[1892]}), .top_right({trees[1893], lumberyards[1893]}), .left({trees[1941], lumberyards[1941]}), .right({trees[1943], lumberyards[1943]}), .bottom_left({trees[1991], lumberyards[1991]}), .bottom({trees[1992], lumberyards[1992]}), .bottom_right({trees[1993], lumberyards[1993]}), .init(2'b01), .state({trees[1942], lumberyards[1942]}));
acre acre_38_43 (.clk(clk), .en(en), .top_left({trees[1892], lumberyards[1892]}), .top({trees[1893], lumberyards[1893]}), .top_right({trees[1894], lumberyards[1894]}), .left({trees[1942], lumberyards[1942]}), .right({trees[1944], lumberyards[1944]}), .bottom_left({trees[1992], lumberyards[1992]}), .bottom({trees[1993], lumberyards[1993]}), .bottom_right({trees[1994], lumberyards[1994]}), .init(2'b00), .state({trees[1943], lumberyards[1943]}));
acre acre_38_44 (.clk(clk), .en(en), .top_left({trees[1893], lumberyards[1893]}), .top({trees[1894], lumberyards[1894]}), .top_right({trees[1895], lumberyards[1895]}), .left({trees[1943], lumberyards[1943]}), .right({trees[1945], lumberyards[1945]}), .bottom_left({trees[1993], lumberyards[1993]}), .bottom({trees[1994], lumberyards[1994]}), .bottom_right({trees[1995], lumberyards[1995]}), .init(2'b00), .state({trees[1944], lumberyards[1944]}));
acre acre_38_45 (.clk(clk), .en(en), .top_left({trees[1894], lumberyards[1894]}), .top({trees[1895], lumberyards[1895]}), .top_right({trees[1896], lumberyards[1896]}), .left({trees[1944], lumberyards[1944]}), .right({trees[1946], lumberyards[1946]}), .bottom_left({trees[1994], lumberyards[1994]}), .bottom({trees[1995], lumberyards[1995]}), .bottom_right({trees[1996], lumberyards[1996]}), .init(2'b10), .state({trees[1945], lumberyards[1945]}));
acre acre_38_46 (.clk(clk), .en(en), .top_left({trees[1895], lumberyards[1895]}), .top({trees[1896], lumberyards[1896]}), .top_right({trees[1897], lumberyards[1897]}), .left({trees[1945], lumberyards[1945]}), .right({trees[1947], lumberyards[1947]}), .bottom_left({trees[1995], lumberyards[1995]}), .bottom({trees[1996], lumberyards[1996]}), .bottom_right({trees[1997], lumberyards[1997]}), .init(2'b10), .state({trees[1946], lumberyards[1946]}));
acre acre_38_47 (.clk(clk), .en(en), .top_left({trees[1896], lumberyards[1896]}), .top({trees[1897], lumberyards[1897]}), .top_right({trees[1898], lumberyards[1898]}), .left({trees[1946], lumberyards[1946]}), .right({trees[1948], lumberyards[1948]}), .bottom_left({trees[1996], lumberyards[1996]}), .bottom({trees[1997], lumberyards[1997]}), .bottom_right({trees[1998], lumberyards[1998]}), .init(2'b00), .state({trees[1947], lumberyards[1947]}));
acre acre_38_48 (.clk(clk), .en(en), .top_left({trees[1897], lumberyards[1897]}), .top({trees[1898], lumberyards[1898]}), .top_right({trees[1899], lumberyards[1899]}), .left({trees[1947], lumberyards[1947]}), .right({trees[1949], lumberyards[1949]}), .bottom_left({trees[1997], lumberyards[1997]}), .bottom({trees[1998], lumberyards[1998]}), .bottom_right({trees[1999], lumberyards[1999]}), .init(2'b00), .state({trees[1948], lumberyards[1948]}));
acre acre_38_49 (.clk(clk), .en(en), .top_left({trees[1898], lumberyards[1898]}), .top({trees[1899], lumberyards[1899]}), .top_right(2'b0), .left({trees[1948], lumberyards[1948]}), .right(2'b0), .bottom_left({trees[1998], lumberyards[1998]}), .bottom({trees[1999], lumberyards[1999]}), .bottom_right(2'b0), .init(2'b00), .state({trees[1949], lumberyards[1949]}));
acre acre_39_0 (.clk(clk), .en(en), .top_left(2'b0), .top({trees[1900], lumberyards[1900]}), .top_right({trees[1901], lumberyards[1901]}), .left(2'b0), .right({trees[1951], lumberyards[1951]}), .bottom_left(2'b0), .bottom({trees[2000], lumberyards[2000]}), .bottom_right({trees[2001], lumberyards[2001]}), .init(2'b00), .state({trees[1950], lumberyards[1950]}));
acre acre_39_1 (.clk(clk), .en(en), .top_left({trees[1900], lumberyards[1900]}), .top({trees[1901], lumberyards[1901]}), .top_right({trees[1902], lumberyards[1902]}), .left({trees[1950], lumberyards[1950]}), .right({trees[1952], lumberyards[1952]}), .bottom_left({trees[2000], lumberyards[2000]}), .bottom({trees[2001], lumberyards[2001]}), .bottom_right({trees[2002], lumberyards[2002]}), .init(2'b00), .state({trees[1951], lumberyards[1951]}));
acre acre_39_2 (.clk(clk), .en(en), .top_left({trees[1901], lumberyards[1901]}), .top({trees[1902], lumberyards[1902]}), .top_right({trees[1903], lumberyards[1903]}), .left({trees[1951], lumberyards[1951]}), .right({trees[1953], lumberyards[1953]}), .bottom_left({trees[2001], lumberyards[2001]}), .bottom({trees[2002], lumberyards[2002]}), .bottom_right({trees[2003], lumberyards[2003]}), .init(2'b00), .state({trees[1952], lumberyards[1952]}));
acre acre_39_3 (.clk(clk), .en(en), .top_left({trees[1902], lumberyards[1902]}), .top({trees[1903], lumberyards[1903]}), .top_right({trees[1904], lumberyards[1904]}), .left({trees[1952], lumberyards[1952]}), .right({trees[1954], lumberyards[1954]}), .bottom_left({trees[2002], lumberyards[2002]}), .bottom({trees[2003], lumberyards[2003]}), .bottom_right({trees[2004], lumberyards[2004]}), .init(2'b10), .state({trees[1953], lumberyards[1953]}));
acre acre_39_4 (.clk(clk), .en(en), .top_left({trees[1903], lumberyards[1903]}), .top({trees[1904], lumberyards[1904]}), .top_right({trees[1905], lumberyards[1905]}), .left({trees[1953], lumberyards[1953]}), .right({trees[1955], lumberyards[1955]}), .bottom_left({trees[2003], lumberyards[2003]}), .bottom({trees[2004], lumberyards[2004]}), .bottom_right({trees[2005], lumberyards[2005]}), .init(2'b10), .state({trees[1954], lumberyards[1954]}));
acre acre_39_5 (.clk(clk), .en(en), .top_left({trees[1904], lumberyards[1904]}), .top({trees[1905], lumberyards[1905]}), .top_right({trees[1906], lumberyards[1906]}), .left({trees[1954], lumberyards[1954]}), .right({trees[1956], lumberyards[1956]}), .bottom_left({trees[2004], lumberyards[2004]}), .bottom({trees[2005], lumberyards[2005]}), .bottom_right({trees[2006], lumberyards[2006]}), .init(2'b01), .state({trees[1955], lumberyards[1955]}));
acre acre_39_6 (.clk(clk), .en(en), .top_left({trees[1905], lumberyards[1905]}), .top({trees[1906], lumberyards[1906]}), .top_right({trees[1907], lumberyards[1907]}), .left({trees[1955], lumberyards[1955]}), .right({trees[1957], lumberyards[1957]}), .bottom_left({trees[2005], lumberyards[2005]}), .bottom({trees[2006], lumberyards[2006]}), .bottom_right({trees[2007], lumberyards[2007]}), .init(2'b10), .state({trees[1956], lumberyards[1956]}));
acre acre_39_7 (.clk(clk), .en(en), .top_left({trees[1906], lumberyards[1906]}), .top({trees[1907], lumberyards[1907]}), .top_right({trees[1908], lumberyards[1908]}), .left({trees[1956], lumberyards[1956]}), .right({trees[1958], lumberyards[1958]}), .bottom_left({trees[2006], lumberyards[2006]}), .bottom({trees[2007], lumberyards[2007]}), .bottom_right({trees[2008], lumberyards[2008]}), .init(2'b00), .state({trees[1957], lumberyards[1957]}));
acre acre_39_8 (.clk(clk), .en(en), .top_left({trees[1907], lumberyards[1907]}), .top({trees[1908], lumberyards[1908]}), .top_right({trees[1909], lumberyards[1909]}), .left({trees[1957], lumberyards[1957]}), .right({trees[1959], lumberyards[1959]}), .bottom_left({trees[2007], lumberyards[2007]}), .bottom({trees[2008], lumberyards[2008]}), .bottom_right({trees[2009], lumberyards[2009]}), .init(2'b00), .state({trees[1958], lumberyards[1958]}));
acre acre_39_9 (.clk(clk), .en(en), .top_left({trees[1908], lumberyards[1908]}), .top({trees[1909], lumberyards[1909]}), .top_right({trees[1910], lumberyards[1910]}), .left({trees[1958], lumberyards[1958]}), .right({trees[1960], lumberyards[1960]}), .bottom_left({trees[2008], lumberyards[2008]}), .bottom({trees[2009], lumberyards[2009]}), .bottom_right({trees[2010], lumberyards[2010]}), .init(2'b00), .state({trees[1959], lumberyards[1959]}));
acre acre_39_10 (.clk(clk), .en(en), .top_left({trees[1909], lumberyards[1909]}), .top({trees[1910], lumberyards[1910]}), .top_right({trees[1911], lumberyards[1911]}), .left({trees[1959], lumberyards[1959]}), .right({trees[1961], lumberyards[1961]}), .bottom_left({trees[2009], lumberyards[2009]}), .bottom({trees[2010], lumberyards[2010]}), .bottom_right({trees[2011], lumberyards[2011]}), .init(2'b10), .state({trees[1960], lumberyards[1960]}));
acre acre_39_11 (.clk(clk), .en(en), .top_left({trees[1910], lumberyards[1910]}), .top({trees[1911], lumberyards[1911]}), .top_right({trees[1912], lumberyards[1912]}), .left({trees[1960], lumberyards[1960]}), .right({trees[1962], lumberyards[1962]}), .bottom_left({trees[2010], lumberyards[2010]}), .bottom({trees[2011], lumberyards[2011]}), .bottom_right({trees[2012], lumberyards[2012]}), .init(2'b00), .state({trees[1961], lumberyards[1961]}));
acre acre_39_12 (.clk(clk), .en(en), .top_left({trees[1911], lumberyards[1911]}), .top({trees[1912], lumberyards[1912]}), .top_right({trees[1913], lumberyards[1913]}), .left({trees[1961], lumberyards[1961]}), .right({trees[1963], lumberyards[1963]}), .bottom_left({trees[2011], lumberyards[2011]}), .bottom({trees[2012], lumberyards[2012]}), .bottom_right({trees[2013], lumberyards[2013]}), .init(2'b01), .state({trees[1962], lumberyards[1962]}));
acre acre_39_13 (.clk(clk), .en(en), .top_left({trees[1912], lumberyards[1912]}), .top({trees[1913], lumberyards[1913]}), .top_right({trees[1914], lumberyards[1914]}), .left({trees[1962], lumberyards[1962]}), .right({trees[1964], lumberyards[1964]}), .bottom_left({trees[2012], lumberyards[2012]}), .bottom({trees[2013], lumberyards[2013]}), .bottom_right({trees[2014], lumberyards[2014]}), .init(2'b00), .state({trees[1963], lumberyards[1963]}));
acre acre_39_14 (.clk(clk), .en(en), .top_left({trees[1913], lumberyards[1913]}), .top({trees[1914], lumberyards[1914]}), .top_right({trees[1915], lumberyards[1915]}), .left({trees[1963], lumberyards[1963]}), .right({trees[1965], lumberyards[1965]}), .bottom_left({trees[2013], lumberyards[2013]}), .bottom({trees[2014], lumberyards[2014]}), .bottom_right({trees[2015], lumberyards[2015]}), .init(2'b00), .state({trees[1964], lumberyards[1964]}));
acre acre_39_15 (.clk(clk), .en(en), .top_left({trees[1914], lumberyards[1914]}), .top({trees[1915], lumberyards[1915]}), .top_right({trees[1916], lumberyards[1916]}), .left({trees[1964], lumberyards[1964]}), .right({trees[1966], lumberyards[1966]}), .bottom_left({trees[2014], lumberyards[2014]}), .bottom({trees[2015], lumberyards[2015]}), .bottom_right({trees[2016], lumberyards[2016]}), .init(2'b10), .state({trees[1965], lumberyards[1965]}));
acre acre_39_16 (.clk(clk), .en(en), .top_left({trees[1915], lumberyards[1915]}), .top({trees[1916], lumberyards[1916]}), .top_right({trees[1917], lumberyards[1917]}), .left({trees[1965], lumberyards[1965]}), .right({trees[1967], lumberyards[1967]}), .bottom_left({trees[2015], lumberyards[2015]}), .bottom({trees[2016], lumberyards[2016]}), .bottom_right({trees[2017], lumberyards[2017]}), .init(2'b00), .state({trees[1966], lumberyards[1966]}));
acre acre_39_17 (.clk(clk), .en(en), .top_left({trees[1916], lumberyards[1916]}), .top({trees[1917], lumberyards[1917]}), .top_right({trees[1918], lumberyards[1918]}), .left({trees[1966], lumberyards[1966]}), .right({trees[1968], lumberyards[1968]}), .bottom_left({trees[2016], lumberyards[2016]}), .bottom({trees[2017], lumberyards[2017]}), .bottom_right({trees[2018], lumberyards[2018]}), .init(2'b01), .state({trees[1967], lumberyards[1967]}));
acre acre_39_18 (.clk(clk), .en(en), .top_left({trees[1917], lumberyards[1917]}), .top({trees[1918], lumberyards[1918]}), .top_right({trees[1919], lumberyards[1919]}), .left({trees[1967], lumberyards[1967]}), .right({trees[1969], lumberyards[1969]}), .bottom_left({trees[2017], lumberyards[2017]}), .bottom({trees[2018], lumberyards[2018]}), .bottom_right({trees[2019], lumberyards[2019]}), .init(2'b00), .state({trees[1968], lumberyards[1968]}));
acre acre_39_19 (.clk(clk), .en(en), .top_left({trees[1918], lumberyards[1918]}), .top({trees[1919], lumberyards[1919]}), .top_right({trees[1920], lumberyards[1920]}), .left({trees[1968], lumberyards[1968]}), .right({trees[1970], lumberyards[1970]}), .bottom_left({trees[2018], lumberyards[2018]}), .bottom({trees[2019], lumberyards[2019]}), .bottom_right({trees[2020], lumberyards[2020]}), .init(2'b00), .state({trees[1969], lumberyards[1969]}));
acre acre_39_20 (.clk(clk), .en(en), .top_left({trees[1919], lumberyards[1919]}), .top({trees[1920], lumberyards[1920]}), .top_right({trees[1921], lumberyards[1921]}), .left({trees[1969], lumberyards[1969]}), .right({trees[1971], lumberyards[1971]}), .bottom_left({trees[2019], lumberyards[2019]}), .bottom({trees[2020], lumberyards[2020]}), .bottom_right({trees[2021], lumberyards[2021]}), .init(2'b00), .state({trees[1970], lumberyards[1970]}));
acre acre_39_21 (.clk(clk), .en(en), .top_left({trees[1920], lumberyards[1920]}), .top({trees[1921], lumberyards[1921]}), .top_right({trees[1922], lumberyards[1922]}), .left({trees[1970], lumberyards[1970]}), .right({trees[1972], lumberyards[1972]}), .bottom_left({trees[2020], lumberyards[2020]}), .bottom({trees[2021], lumberyards[2021]}), .bottom_right({trees[2022], lumberyards[2022]}), .init(2'b00), .state({trees[1971], lumberyards[1971]}));
acre acre_39_22 (.clk(clk), .en(en), .top_left({trees[1921], lumberyards[1921]}), .top({trees[1922], lumberyards[1922]}), .top_right({trees[1923], lumberyards[1923]}), .left({trees[1971], lumberyards[1971]}), .right({trees[1973], lumberyards[1973]}), .bottom_left({trees[2021], lumberyards[2021]}), .bottom({trees[2022], lumberyards[2022]}), .bottom_right({trees[2023], lumberyards[2023]}), .init(2'b00), .state({trees[1972], lumberyards[1972]}));
acre acre_39_23 (.clk(clk), .en(en), .top_left({trees[1922], lumberyards[1922]}), .top({trees[1923], lumberyards[1923]}), .top_right({trees[1924], lumberyards[1924]}), .left({trees[1972], lumberyards[1972]}), .right({trees[1974], lumberyards[1974]}), .bottom_left({trees[2022], lumberyards[2022]}), .bottom({trees[2023], lumberyards[2023]}), .bottom_right({trees[2024], lumberyards[2024]}), .init(2'b01), .state({trees[1973], lumberyards[1973]}));
acre acre_39_24 (.clk(clk), .en(en), .top_left({trees[1923], lumberyards[1923]}), .top({trees[1924], lumberyards[1924]}), .top_right({trees[1925], lumberyards[1925]}), .left({trees[1973], lumberyards[1973]}), .right({trees[1975], lumberyards[1975]}), .bottom_left({trees[2023], lumberyards[2023]}), .bottom({trees[2024], lumberyards[2024]}), .bottom_right({trees[2025], lumberyards[2025]}), .init(2'b00), .state({trees[1974], lumberyards[1974]}));
acre acre_39_25 (.clk(clk), .en(en), .top_left({trees[1924], lumberyards[1924]}), .top({trees[1925], lumberyards[1925]}), .top_right({trees[1926], lumberyards[1926]}), .left({trees[1974], lumberyards[1974]}), .right({trees[1976], lumberyards[1976]}), .bottom_left({trees[2024], lumberyards[2024]}), .bottom({trees[2025], lumberyards[2025]}), .bottom_right({trees[2026], lumberyards[2026]}), .init(2'b00), .state({trees[1975], lumberyards[1975]}));
acre acre_39_26 (.clk(clk), .en(en), .top_left({trees[1925], lumberyards[1925]}), .top({trees[1926], lumberyards[1926]}), .top_right({trees[1927], lumberyards[1927]}), .left({trees[1975], lumberyards[1975]}), .right({trees[1977], lumberyards[1977]}), .bottom_left({trees[2025], lumberyards[2025]}), .bottom({trees[2026], lumberyards[2026]}), .bottom_right({trees[2027], lumberyards[2027]}), .init(2'b00), .state({trees[1976], lumberyards[1976]}));
acre acre_39_27 (.clk(clk), .en(en), .top_left({trees[1926], lumberyards[1926]}), .top({trees[1927], lumberyards[1927]}), .top_right({trees[1928], lumberyards[1928]}), .left({trees[1976], lumberyards[1976]}), .right({trees[1978], lumberyards[1978]}), .bottom_left({trees[2026], lumberyards[2026]}), .bottom({trees[2027], lumberyards[2027]}), .bottom_right({trees[2028], lumberyards[2028]}), .init(2'b00), .state({trees[1977], lumberyards[1977]}));
acre acre_39_28 (.clk(clk), .en(en), .top_left({trees[1927], lumberyards[1927]}), .top({trees[1928], lumberyards[1928]}), .top_right({trees[1929], lumberyards[1929]}), .left({trees[1977], lumberyards[1977]}), .right({trees[1979], lumberyards[1979]}), .bottom_left({trees[2027], lumberyards[2027]}), .bottom({trees[2028], lumberyards[2028]}), .bottom_right({trees[2029], lumberyards[2029]}), .init(2'b00), .state({trees[1978], lumberyards[1978]}));
acre acre_39_29 (.clk(clk), .en(en), .top_left({trees[1928], lumberyards[1928]}), .top({trees[1929], lumberyards[1929]}), .top_right({trees[1930], lumberyards[1930]}), .left({trees[1978], lumberyards[1978]}), .right({trees[1980], lumberyards[1980]}), .bottom_left({trees[2028], lumberyards[2028]}), .bottom({trees[2029], lumberyards[2029]}), .bottom_right({trees[2030], lumberyards[2030]}), .init(2'b01), .state({trees[1979], lumberyards[1979]}));
acre acre_39_30 (.clk(clk), .en(en), .top_left({trees[1929], lumberyards[1929]}), .top({trees[1930], lumberyards[1930]}), .top_right({trees[1931], lumberyards[1931]}), .left({trees[1979], lumberyards[1979]}), .right({trees[1981], lumberyards[1981]}), .bottom_left({trees[2029], lumberyards[2029]}), .bottom({trees[2030], lumberyards[2030]}), .bottom_right({trees[2031], lumberyards[2031]}), .init(2'b00), .state({trees[1980], lumberyards[1980]}));
acre acre_39_31 (.clk(clk), .en(en), .top_left({trees[1930], lumberyards[1930]}), .top({trees[1931], lumberyards[1931]}), .top_right({trees[1932], lumberyards[1932]}), .left({trees[1980], lumberyards[1980]}), .right({trees[1982], lumberyards[1982]}), .bottom_left({trees[2030], lumberyards[2030]}), .bottom({trees[2031], lumberyards[2031]}), .bottom_right({trees[2032], lumberyards[2032]}), .init(2'b01), .state({trees[1981], lumberyards[1981]}));
acre acre_39_32 (.clk(clk), .en(en), .top_left({trees[1931], lumberyards[1931]}), .top({trees[1932], lumberyards[1932]}), .top_right({trees[1933], lumberyards[1933]}), .left({trees[1981], lumberyards[1981]}), .right({trees[1983], lumberyards[1983]}), .bottom_left({trees[2031], lumberyards[2031]}), .bottom({trees[2032], lumberyards[2032]}), .bottom_right({trees[2033], lumberyards[2033]}), .init(2'b00), .state({trees[1982], lumberyards[1982]}));
acre acre_39_33 (.clk(clk), .en(en), .top_left({trees[1932], lumberyards[1932]}), .top({trees[1933], lumberyards[1933]}), .top_right({trees[1934], lumberyards[1934]}), .left({trees[1982], lumberyards[1982]}), .right({trees[1984], lumberyards[1984]}), .bottom_left({trees[2032], lumberyards[2032]}), .bottom({trees[2033], lumberyards[2033]}), .bottom_right({trees[2034], lumberyards[2034]}), .init(2'b01), .state({trees[1983], lumberyards[1983]}));
acre acre_39_34 (.clk(clk), .en(en), .top_left({trees[1933], lumberyards[1933]}), .top({trees[1934], lumberyards[1934]}), .top_right({trees[1935], lumberyards[1935]}), .left({trees[1983], lumberyards[1983]}), .right({trees[1985], lumberyards[1985]}), .bottom_left({trees[2033], lumberyards[2033]}), .bottom({trees[2034], lumberyards[2034]}), .bottom_right({trees[2035], lumberyards[2035]}), .init(2'b00), .state({trees[1984], lumberyards[1984]}));
acre acre_39_35 (.clk(clk), .en(en), .top_left({trees[1934], lumberyards[1934]}), .top({trees[1935], lumberyards[1935]}), .top_right({trees[1936], lumberyards[1936]}), .left({trees[1984], lumberyards[1984]}), .right({trees[1986], lumberyards[1986]}), .bottom_left({trees[2034], lumberyards[2034]}), .bottom({trees[2035], lumberyards[2035]}), .bottom_right({trees[2036], lumberyards[2036]}), .init(2'b01), .state({trees[1985], lumberyards[1985]}));
acre acre_39_36 (.clk(clk), .en(en), .top_left({trees[1935], lumberyards[1935]}), .top({trees[1936], lumberyards[1936]}), .top_right({trees[1937], lumberyards[1937]}), .left({trees[1985], lumberyards[1985]}), .right({trees[1987], lumberyards[1987]}), .bottom_left({trees[2035], lumberyards[2035]}), .bottom({trees[2036], lumberyards[2036]}), .bottom_right({trees[2037], lumberyards[2037]}), .init(2'b01), .state({trees[1986], lumberyards[1986]}));
acre acre_39_37 (.clk(clk), .en(en), .top_left({trees[1936], lumberyards[1936]}), .top({trees[1937], lumberyards[1937]}), .top_right({trees[1938], lumberyards[1938]}), .left({trees[1986], lumberyards[1986]}), .right({trees[1988], lumberyards[1988]}), .bottom_left({trees[2036], lumberyards[2036]}), .bottom({trees[2037], lumberyards[2037]}), .bottom_right({trees[2038], lumberyards[2038]}), .init(2'b00), .state({trees[1987], lumberyards[1987]}));
acre acre_39_38 (.clk(clk), .en(en), .top_left({trees[1937], lumberyards[1937]}), .top({trees[1938], lumberyards[1938]}), .top_right({trees[1939], lumberyards[1939]}), .left({trees[1987], lumberyards[1987]}), .right({trees[1989], lumberyards[1989]}), .bottom_left({trees[2037], lumberyards[2037]}), .bottom({trees[2038], lumberyards[2038]}), .bottom_right({trees[2039], lumberyards[2039]}), .init(2'b00), .state({trees[1988], lumberyards[1988]}));
acre acre_39_39 (.clk(clk), .en(en), .top_left({trees[1938], lumberyards[1938]}), .top({trees[1939], lumberyards[1939]}), .top_right({trees[1940], lumberyards[1940]}), .left({trees[1988], lumberyards[1988]}), .right({trees[1990], lumberyards[1990]}), .bottom_left({trees[2038], lumberyards[2038]}), .bottom({trees[2039], lumberyards[2039]}), .bottom_right({trees[2040], lumberyards[2040]}), .init(2'b01), .state({trees[1989], lumberyards[1989]}));
acre acre_39_40 (.clk(clk), .en(en), .top_left({trees[1939], lumberyards[1939]}), .top({trees[1940], lumberyards[1940]}), .top_right({trees[1941], lumberyards[1941]}), .left({trees[1989], lumberyards[1989]}), .right({trees[1991], lumberyards[1991]}), .bottom_left({trees[2039], lumberyards[2039]}), .bottom({trees[2040], lumberyards[2040]}), .bottom_right({trees[2041], lumberyards[2041]}), .init(2'b00), .state({trees[1990], lumberyards[1990]}));
acre acre_39_41 (.clk(clk), .en(en), .top_left({trees[1940], lumberyards[1940]}), .top({trees[1941], lumberyards[1941]}), .top_right({trees[1942], lumberyards[1942]}), .left({trees[1990], lumberyards[1990]}), .right({trees[1992], lumberyards[1992]}), .bottom_left({trees[2040], lumberyards[2040]}), .bottom({trees[2041], lumberyards[2041]}), .bottom_right({trees[2042], lumberyards[2042]}), .init(2'b00), .state({trees[1991], lumberyards[1991]}));
acre acre_39_42 (.clk(clk), .en(en), .top_left({trees[1941], lumberyards[1941]}), .top({trees[1942], lumberyards[1942]}), .top_right({trees[1943], lumberyards[1943]}), .left({trees[1991], lumberyards[1991]}), .right({trees[1993], lumberyards[1993]}), .bottom_left({trees[2041], lumberyards[2041]}), .bottom({trees[2042], lumberyards[2042]}), .bottom_right({trees[2043], lumberyards[2043]}), .init(2'b00), .state({trees[1992], lumberyards[1992]}));
acre acre_39_43 (.clk(clk), .en(en), .top_left({trees[1942], lumberyards[1942]}), .top({trees[1943], lumberyards[1943]}), .top_right({trees[1944], lumberyards[1944]}), .left({trees[1992], lumberyards[1992]}), .right({trees[1994], lumberyards[1994]}), .bottom_left({trees[2042], lumberyards[2042]}), .bottom({trees[2043], lumberyards[2043]}), .bottom_right({trees[2044], lumberyards[2044]}), .init(2'b00), .state({trees[1993], lumberyards[1993]}));
acre acre_39_44 (.clk(clk), .en(en), .top_left({trees[1943], lumberyards[1943]}), .top({trees[1944], lumberyards[1944]}), .top_right({trees[1945], lumberyards[1945]}), .left({trees[1993], lumberyards[1993]}), .right({trees[1995], lumberyards[1995]}), .bottom_left({trees[2043], lumberyards[2043]}), .bottom({trees[2044], lumberyards[2044]}), .bottom_right({trees[2045], lumberyards[2045]}), .init(2'b10), .state({trees[1994], lumberyards[1994]}));
acre acre_39_45 (.clk(clk), .en(en), .top_left({trees[1944], lumberyards[1944]}), .top({trees[1945], lumberyards[1945]}), .top_right({trees[1946], lumberyards[1946]}), .left({trees[1994], lumberyards[1994]}), .right({trees[1996], lumberyards[1996]}), .bottom_left({trees[2044], lumberyards[2044]}), .bottom({trees[2045], lumberyards[2045]}), .bottom_right({trees[2046], lumberyards[2046]}), .init(2'b00), .state({trees[1995], lumberyards[1995]}));
acre acre_39_46 (.clk(clk), .en(en), .top_left({trees[1945], lumberyards[1945]}), .top({trees[1946], lumberyards[1946]}), .top_right({trees[1947], lumberyards[1947]}), .left({trees[1995], lumberyards[1995]}), .right({trees[1997], lumberyards[1997]}), .bottom_left({trees[2045], lumberyards[2045]}), .bottom({trees[2046], lumberyards[2046]}), .bottom_right({trees[2047], lumberyards[2047]}), .init(2'b00), .state({trees[1996], lumberyards[1996]}));
acre acre_39_47 (.clk(clk), .en(en), .top_left({trees[1946], lumberyards[1946]}), .top({trees[1947], lumberyards[1947]}), .top_right({trees[1948], lumberyards[1948]}), .left({trees[1996], lumberyards[1996]}), .right({trees[1998], lumberyards[1998]}), .bottom_left({trees[2046], lumberyards[2046]}), .bottom({trees[2047], lumberyards[2047]}), .bottom_right({trees[2048], lumberyards[2048]}), .init(2'b01), .state({trees[1997], lumberyards[1997]}));
acre acre_39_48 (.clk(clk), .en(en), .top_left({trees[1947], lumberyards[1947]}), .top({trees[1948], lumberyards[1948]}), .top_right({trees[1949], lumberyards[1949]}), .left({trees[1997], lumberyards[1997]}), .right({trees[1999], lumberyards[1999]}), .bottom_left({trees[2047], lumberyards[2047]}), .bottom({trees[2048], lumberyards[2048]}), .bottom_right({trees[2049], lumberyards[2049]}), .init(2'b10), .state({trees[1998], lumberyards[1998]}));
acre acre_39_49 (.clk(clk), .en(en), .top_left({trees[1948], lumberyards[1948]}), .top({trees[1949], lumberyards[1949]}), .top_right(2'b0), .left({trees[1998], lumberyards[1998]}), .right(2'b0), .bottom_left({trees[2048], lumberyards[2048]}), .bottom({trees[2049], lumberyards[2049]}), .bottom_right(2'b0), .init(2'b00), .state({trees[1999], lumberyards[1999]}));
acre acre_40_0 (.clk(clk), .en(en), .top_left(2'b0), .top({trees[1950], lumberyards[1950]}), .top_right({trees[1951], lumberyards[1951]}), .left(2'b0), .right({trees[2001], lumberyards[2001]}), .bottom_left(2'b0), .bottom({trees[2050], lumberyards[2050]}), .bottom_right({trees[2051], lumberyards[2051]}), .init(2'b01), .state({trees[2000], lumberyards[2000]}));
acre acre_40_1 (.clk(clk), .en(en), .top_left({trees[1950], lumberyards[1950]}), .top({trees[1951], lumberyards[1951]}), .top_right({trees[1952], lumberyards[1952]}), .left({trees[2000], lumberyards[2000]}), .right({trees[2002], lumberyards[2002]}), .bottom_left({trees[2050], lumberyards[2050]}), .bottom({trees[2051], lumberyards[2051]}), .bottom_right({trees[2052], lumberyards[2052]}), .init(2'b00), .state({trees[2001], lumberyards[2001]}));
acre acre_40_2 (.clk(clk), .en(en), .top_left({trees[1951], lumberyards[1951]}), .top({trees[1952], lumberyards[1952]}), .top_right({trees[1953], lumberyards[1953]}), .left({trees[2001], lumberyards[2001]}), .right({trees[2003], lumberyards[2003]}), .bottom_left({trees[2051], lumberyards[2051]}), .bottom({trees[2052], lumberyards[2052]}), .bottom_right({trees[2053], lumberyards[2053]}), .init(2'b01), .state({trees[2002], lumberyards[2002]}));
acre acre_40_3 (.clk(clk), .en(en), .top_left({trees[1952], lumberyards[1952]}), .top({trees[1953], lumberyards[1953]}), .top_right({trees[1954], lumberyards[1954]}), .left({trees[2002], lumberyards[2002]}), .right({trees[2004], lumberyards[2004]}), .bottom_left({trees[2052], lumberyards[2052]}), .bottom({trees[2053], lumberyards[2053]}), .bottom_right({trees[2054], lumberyards[2054]}), .init(2'b01), .state({trees[2003], lumberyards[2003]}));
acre acre_40_4 (.clk(clk), .en(en), .top_left({trees[1953], lumberyards[1953]}), .top({trees[1954], lumberyards[1954]}), .top_right({trees[1955], lumberyards[1955]}), .left({trees[2003], lumberyards[2003]}), .right({trees[2005], lumberyards[2005]}), .bottom_left({trees[2053], lumberyards[2053]}), .bottom({trees[2054], lumberyards[2054]}), .bottom_right({trees[2055], lumberyards[2055]}), .init(2'b10), .state({trees[2004], lumberyards[2004]}));
acre acre_40_5 (.clk(clk), .en(en), .top_left({trees[1954], lumberyards[1954]}), .top({trees[1955], lumberyards[1955]}), .top_right({trees[1956], lumberyards[1956]}), .left({trees[2004], lumberyards[2004]}), .right({trees[2006], lumberyards[2006]}), .bottom_left({trees[2054], lumberyards[2054]}), .bottom({trees[2055], lumberyards[2055]}), .bottom_right({trees[2056], lumberyards[2056]}), .init(2'b00), .state({trees[2005], lumberyards[2005]}));
acre acre_40_6 (.clk(clk), .en(en), .top_left({trees[1955], lumberyards[1955]}), .top({trees[1956], lumberyards[1956]}), .top_right({trees[1957], lumberyards[1957]}), .left({trees[2005], lumberyards[2005]}), .right({trees[2007], lumberyards[2007]}), .bottom_left({trees[2055], lumberyards[2055]}), .bottom({trees[2056], lumberyards[2056]}), .bottom_right({trees[2057], lumberyards[2057]}), .init(2'b00), .state({trees[2006], lumberyards[2006]}));
acre acre_40_7 (.clk(clk), .en(en), .top_left({trees[1956], lumberyards[1956]}), .top({trees[1957], lumberyards[1957]}), .top_right({trees[1958], lumberyards[1958]}), .left({trees[2006], lumberyards[2006]}), .right({trees[2008], lumberyards[2008]}), .bottom_left({trees[2056], lumberyards[2056]}), .bottom({trees[2057], lumberyards[2057]}), .bottom_right({trees[2058], lumberyards[2058]}), .init(2'b00), .state({trees[2007], lumberyards[2007]}));
acre acre_40_8 (.clk(clk), .en(en), .top_left({trees[1957], lumberyards[1957]}), .top({trees[1958], lumberyards[1958]}), .top_right({trees[1959], lumberyards[1959]}), .left({trees[2007], lumberyards[2007]}), .right({trees[2009], lumberyards[2009]}), .bottom_left({trees[2057], lumberyards[2057]}), .bottom({trees[2058], lumberyards[2058]}), .bottom_right({trees[2059], lumberyards[2059]}), .init(2'b00), .state({trees[2008], lumberyards[2008]}));
acre acre_40_9 (.clk(clk), .en(en), .top_left({trees[1958], lumberyards[1958]}), .top({trees[1959], lumberyards[1959]}), .top_right({trees[1960], lumberyards[1960]}), .left({trees[2008], lumberyards[2008]}), .right({trees[2010], lumberyards[2010]}), .bottom_left({trees[2058], lumberyards[2058]}), .bottom({trees[2059], lumberyards[2059]}), .bottom_right({trees[2060], lumberyards[2060]}), .init(2'b10), .state({trees[2009], lumberyards[2009]}));
acre acre_40_10 (.clk(clk), .en(en), .top_left({trees[1959], lumberyards[1959]}), .top({trees[1960], lumberyards[1960]}), .top_right({trees[1961], lumberyards[1961]}), .left({trees[2009], lumberyards[2009]}), .right({trees[2011], lumberyards[2011]}), .bottom_left({trees[2059], lumberyards[2059]}), .bottom({trees[2060], lumberyards[2060]}), .bottom_right({trees[2061], lumberyards[2061]}), .init(2'b00), .state({trees[2010], lumberyards[2010]}));
acre acre_40_11 (.clk(clk), .en(en), .top_left({trees[1960], lumberyards[1960]}), .top({trees[1961], lumberyards[1961]}), .top_right({trees[1962], lumberyards[1962]}), .left({trees[2010], lumberyards[2010]}), .right({trees[2012], lumberyards[2012]}), .bottom_left({trees[2060], lumberyards[2060]}), .bottom({trees[2061], lumberyards[2061]}), .bottom_right({trees[2062], lumberyards[2062]}), .init(2'b10), .state({trees[2011], lumberyards[2011]}));
acre acre_40_12 (.clk(clk), .en(en), .top_left({trees[1961], lumberyards[1961]}), .top({trees[1962], lumberyards[1962]}), .top_right({trees[1963], lumberyards[1963]}), .left({trees[2011], lumberyards[2011]}), .right({trees[2013], lumberyards[2013]}), .bottom_left({trees[2061], lumberyards[2061]}), .bottom({trees[2062], lumberyards[2062]}), .bottom_right({trees[2063], lumberyards[2063]}), .init(2'b10), .state({trees[2012], lumberyards[2012]}));
acre acre_40_13 (.clk(clk), .en(en), .top_left({trees[1962], lumberyards[1962]}), .top({trees[1963], lumberyards[1963]}), .top_right({trees[1964], lumberyards[1964]}), .left({trees[2012], lumberyards[2012]}), .right({trees[2014], lumberyards[2014]}), .bottom_left({trees[2062], lumberyards[2062]}), .bottom({trees[2063], lumberyards[2063]}), .bottom_right({trees[2064], lumberyards[2064]}), .init(2'b00), .state({trees[2013], lumberyards[2013]}));
acre acre_40_14 (.clk(clk), .en(en), .top_left({trees[1963], lumberyards[1963]}), .top({trees[1964], lumberyards[1964]}), .top_right({trees[1965], lumberyards[1965]}), .left({trees[2013], lumberyards[2013]}), .right({trees[2015], lumberyards[2015]}), .bottom_left({trees[2063], lumberyards[2063]}), .bottom({trees[2064], lumberyards[2064]}), .bottom_right({trees[2065], lumberyards[2065]}), .init(2'b10), .state({trees[2014], lumberyards[2014]}));
acre acre_40_15 (.clk(clk), .en(en), .top_left({trees[1964], lumberyards[1964]}), .top({trees[1965], lumberyards[1965]}), .top_right({trees[1966], lumberyards[1966]}), .left({trees[2014], lumberyards[2014]}), .right({trees[2016], lumberyards[2016]}), .bottom_left({trees[2064], lumberyards[2064]}), .bottom({trees[2065], lumberyards[2065]}), .bottom_right({trees[2066], lumberyards[2066]}), .init(2'b00), .state({trees[2015], lumberyards[2015]}));
acre acre_40_16 (.clk(clk), .en(en), .top_left({trees[1965], lumberyards[1965]}), .top({trees[1966], lumberyards[1966]}), .top_right({trees[1967], lumberyards[1967]}), .left({trees[2015], lumberyards[2015]}), .right({trees[2017], lumberyards[2017]}), .bottom_left({trees[2065], lumberyards[2065]}), .bottom({trees[2066], lumberyards[2066]}), .bottom_right({trees[2067], lumberyards[2067]}), .init(2'b00), .state({trees[2016], lumberyards[2016]}));
acre acre_40_17 (.clk(clk), .en(en), .top_left({trees[1966], lumberyards[1966]}), .top({trees[1967], lumberyards[1967]}), .top_right({trees[1968], lumberyards[1968]}), .left({trees[2016], lumberyards[2016]}), .right({trees[2018], lumberyards[2018]}), .bottom_left({trees[2066], lumberyards[2066]}), .bottom({trees[2067], lumberyards[2067]}), .bottom_right({trees[2068], lumberyards[2068]}), .init(2'b10), .state({trees[2017], lumberyards[2017]}));
acre acre_40_18 (.clk(clk), .en(en), .top_left({trees[1967], lumberyards[1967]}), .top({trees[1968], lumberyards[1968]}), .top_right({trees[1969], lumberyards[1969]}), .left({trees[2017], lumberyards[2017]}), .right({trees[2019], lumberyards[2019]}), .bottom_left({trees[2067], lumberyards[2067]}), .bottom({trees[2068], lumberyards[2068]}), .bottom_right({trees[2069], lumberyards[2069]}), .init(2'b00), .state({trees[2018], lumberyards[2018]}));
acre acre_40_19 (.clk(clk), .en(en), .top_left({trees[1968], lumberyards[1968]}), .top({trees[1969], lumberyards[1969]}), .top_right({trees[1970], lumberyards[1970]}), .left({trees[2018], lumberyards[2018]}), .right({trees[2020], lumberyards[2020]}), .bottom_left({trees[2068], lumberyards[2068]}), .bottom({trees[2069], lumberyards[2069]}), .bottom_right({trees[2070], lumberyards[2070]}), .init(2'b00), .state({trees[2019], lumberyards[2019]}));
acre acre_40_20 (.clk(clk), .en(en), .top_left({trees[1969], lumberyards[1969]}), .top({trees[1970], lumberyards[1970]}), .top_right({trees[1971], lumberyards[1971]}), .left({trees[2019], lumberyards[2019]}), .right({trees[2021], lumberyards[2021]}), .bottom_left({trees[2069], lumberyards[2069]}), .bottom({trees[2070], lumberyards[2070]}), .bottom_right({trees[2071], lumberyards[2071]}), .init(2'b01), .state({trees[2020], lumberyards[2020]}));
acre acre_40_21 (.clk(clk), .en(en), .top_left({trees[1970], lumberyards[1970]}), .top({trees[1971], lumberyards[1971]}), .top_right({trees[1972], lumberyards[1972]}), .left({trees[2020], lumberyards[2020]}), .right({trees[2022], lumberyards[2022]}), .bottom_left({trees[2070], lumberyards[2070]}), .bottom({trees[2071], lumberyards[2071]}), .bottom_right({trees[2072], lumberyards[2072]}), .init(2'b00), .state({trees[2021], lumberyards[2021]}));
acre acre_40_22 (.clk(clk), .en(en), .top_left({trees[1971], lumberyards[1971]}), .top({trees[1972], lumberyards[1972]}), .top_right({trees[1973], lumberyards[1973]}), .left({trees[2021], lumberyards[2021]}), .right({trees[2023], lumberyards[2023]}), .bottom_left({trees[2071], lumberyards[2071]}), .bottom({trees[2072], lumberyards[2072]}), .bottom_right({trees[2073], lumberyards[2073]}), .init(2'b00), .state({trees[2022], lumberyards[2022]}));
acre acre_40_23 (.clk(clk), .en(en), .top_left({trees[1972], lumberyards[1972]}), .top({trees[1973], lumberyards[1973]}), .top_right({trees[1974], lumberyards[1974]}), .left({trees[2022], lumberyards[2022]}), .right({trees[2024], lumberyards[2024]}), .bottom_left({trees[2072], lumberyards[2072]}), .bottom({trees[2073], lumberyards[2073]}), .bottom_right({trees[2074], lumberyards[2074]}), .init(2'b00), .state({trees[2023], lumberyards[2023]}));
acre acre_40_24 (.clk(clk), .en(en), .top_left({trees[1973], lumberyards[1973]}), .top({trees[1974], lumberyards[1974]}), .top_right({trees[1975], lumberyards[1975]}), .left({trees[2023], lumberyards[2023]}), .right({trees[2025], lumberyards[2025]}), .bottom_left({trees[2073], lumberyards[2073]}), .bottom({trees[2074], lumberyards[2074]}), .bottom_right({trees[2075], lumberyards[2075]}), .init(2'b00), .state({trees[2024], lumberyards[2024]}));
acre acre_40_25 (.clk(clk), .en(en), .top_left({trees[1974], lumberyards[1974]}), .top({trees[1975], lumberyards[1975]}), .top_right({trees[1976], lumberyards[1976]}), .left({trees[2024], lumberyards[2024]}), .right({trees[2026], lumberyards[2026]}), .bottom_left({trees[2074], lumberyards[2074]}), .bottom({trees[2075], lumberyards[2075]}), .bottom_right({trees[2076], lumberyards[2076]}), .init(2'b00), .state({trees[2025], lumberyards[2025]}));
acre acre_40_26 (.clk(clk), .en(en), .top_left({trees[1975], lumberyards[1975]}), .top({trees[1976], lumberyards[1976]}), .top_right({trees[1977], lumberyards[1977]}), .left({trees[2025], lumberyards[2025]}), .right({trees[2027], lumberyards[2027]}), .bottom_left({trees[2075], lumberyards[2075]}), .bottom({trees[2076], lumberyards[2076]}), .bottom_right({trees[2077], lumberyards[2077]}), .init(2'b00), .state({trees[2026], lumberyards[2026]}));
acre acre_40_27 (.clk(clk), .en(en), .top_left({trees[1976], lumberyards[1976]}), .top({trees[1977], lumberyards[1977]}), .top_right({trees[1978], lumberyards[1978]}), .left({trees[2026], lumberyards[2026]}), .right({trees[2028], lumberyards[2028]}), .bottom_left({trees[2076], lumberyards[2076]}), .bottom({trees[2077], lumberyards[2077]}), .bottom_right({trees[2078], lumberyards[2078]}), .init(2'b01), .state({trees[2027], lumberyards[2027]}));
acre acre_40_28 (.clk(clk), .en(en), .top_left({trees[1977], lumberyards[1977]}), .top({trees[1978], lumberyards[1978]}), .top_right({trees[1979], lumberyards[1979]}), .left({trees[2027], lumberyards[2027]}), .right({trees[2029], lumberyards[2029]}), .bottom_left({trees[2077], lumberyards[2077]}), .bottom({trees[2078], lumberyards[2078]}), .bottom_right({trees[2079], lumberyards[2079]}), .init(2'b00), .state({trees[2028], lumberyards[2028]}));
acre acre_40_29 (.clk(clk), .en(en), .top_left({trees[1978], lumberyards[1978]}), .top({trees[1979], lumberyards[1979]}), .top_right({trees[1980], lumberyards[1980]}), .left({trees[2028], lumberyards[2028]}), .right({trees[2030], lumberyards[2030]}), .bottom_left({trees[2078], lumberyards[2078]}), .bottom({trees[2079], lumberyards[2079]}), .bottom_right({trees[2080], lumberyards[2080]}), .init(2'b00), .state({trees[2029], lumberyards[2029]}));
acre acre_40_30 (.clk(clk), .en(en), .top_left({trees[1979], lumberyards[1979]}), .top({trees[1980], lumberyards[1980]}), .top_right({trees[1981], lumberyards[1981]}), .left({trees[2029], lumberyards[2029]}), .right({trees[2031], lumberyards[2031]}), .bottom_left({trees[2079], lumberyards[2079]}), .bottom({trees[2080], lumberyards[2080]}), .bottom_right({trees[2081], lumberyards[2081]}), .init(2'b00), .state({trees[2030], lumberyards[2030]}));
acre acre_40_31 (.clk(clk), .en(en), .top_left({trees[1980], lumberyards[1980]}), .top({trees[1981], lumberyards[1981]}), .top_right({trees[1982], lumberyards[1982]}), .left({trees[2030], lumberyards[2030]}), .right({trees[2032], lumberyards[2032]}), .bottom_left({trees[2080], lumberyards[2080]}), .bottom({trees[2081], lumberyards[2081]}), .bottom_right({trees[2082], lumberyards[2082]}), .init(2'b00), .state({trees[2031], lumberyards[2031]}));
acre acre_40_32 (.clk(clk), .en(en), .top_left({trees[1981], lumberyards[1981]}), .top({trees[1982], lumberyards[1982]}), .top_right({trees[1983], lumberyards[1983]}), .left({trees[2031], lumberyards[2031]}), .right({trees[2033], lumberyards[2033]}), .bottom_left({trees[2081], lumberyards[2081]}), .bottom({trees[2082], lumberyards[2082]}), .bottom_right({trees[2083], lumberyards[2083]}), .init(2'b10), .state({trees[2032], lumberyards[2032]}));
acre acre_40_33 (.clk(clk), .en(en), .top_left({trees[1982], lumberyards[1982]}), .top({trees[1983], lumberyards[1983]}), .top_right({trees[1984], lumberyards[1984]}), .left({trees[2032], lumberyards[2032]}), .right({trees[2034], lumberyards[2034]}), .bottom_left({trees[2082], lumberyards[2082]}), .bottom({trees[2083], lumberyards[2083]}), .bottom_right({trees[2084], lumberyards[2084]}), .init(2'b10), .state({trees[2033], lumberyards[2033]}));
acre acre_40_34 (.clk(clk), .en(en), .top_left({trees[1983], lumberyards[1983]}), .top({trees[1984], lumberyards[1984]}), .top_right({trees[1985], lumberyards[1985]}), .left({trees[2033], lumberyards[2033]}), .right({trees[2035], lumberyards[2035]}), .bottom_left({trees[2083], lumberyards[2083]}), .bottom({trees[2084], lumberyards[2084]}), .bottom_right({trees[2085], lumberyards[2085]}), .init(2'b00), .state({trees[2034], lumberyards[2034]}));
acre acre_40_35 (.clk(clk), .en(en), .top_left({trees[1984], lumberyards[1984]}), .top({trees[1985], lumberyards[1985]}), .top_right({trees[1986], lumberyards[1986]}), .left({trees[2034], lumberyards[2034]}), .right({trees[2036], lumberyards[2036]}), .bottom_left({trees[2084], lumberyards[2084]}), .bottom({trees[2085], lumberyards[2085]}), .bottom_right({trees[2086], lumberyards[2086]}), .init(2'b01), .state({trees[2035], lumberyards[2035]}));
acre acre_40_36 (.clk(clk), .en(en), .top_left({trees[1985], lumberyards[1985]}), .top({trees[1986], lumberyards[1986]}), .top_right({trees[1987], lumberyards[1987]}), .left({trees[2035], lumberyards[2035]}), .right({trees[2037], lumberyards[2037]}), .bottom_left({trees[2085], lumberyards[2085]}), .bottom({trees[2086], lumberyards[2086]}), .bottom_right({trees[2087], lumberyards[2087]}), .init(2'b00), .state({trees[2036], lumberyards[2036]}));
acre acre_40_37 (.clk(clk), .en(en), .top_left({trees[1986], lumberyards[1986]}), .top({trees[1987], lumberyards[1987]}), .top_right({trees[1988], lumberyards[1988]}), .left({trees[2036], lumberyards[2036]}), .right({trees[2038], lumberyards[2038]}), .bottom_left({trees[2086], lumberyards[2086]}), .bottom({trees[2087], lumberyards[2087]}), .bottom_right({trees[2088], lumberyards[2088]}), .init(2'b00), .state({trees[2037], lumberyards[2037]}));
acre acre_40_38 (.clk(clk), .en(en), .top_left({trees[1987], lumberyards[1987]}), .top({trees[1988], lumberyards[1988]}), .top_right({trees[1989], lumberyards[1989]}), .left({trees[2037], lumberyards[2037]}), .right({trees[2039], lumberyards[2039]}), .bottom_left({trees[2087], lumberyards[2087]}), .bottom({trees[2088], lumberyards[2088]}), .bottom_right({trees[2089], lumberyards[2089]}), .init(2'b01), .state({trees[2038], lumberyards[2038]}));
acre acre_40_39 (.clk(clk), .en(en), .top_left({trees[1988], lumberyards[1988]}), .top({trees[1989], lumberyards[1989]}), .top_right({trees[1990], lumberyards[1990]}), .left({trees[2038], lumberyards[2038]}), .right({trees[2040], lumberyards[2040]}), .bottom_left({trees[2088], lumberyards[2088]}), .bottom({trees[2089], lumberyards[2089]}), .bottom_right({trees[2090], lumberyards[2090]}), .init(2'b01), .state({trees[2039], lumberyards[2039]}));
acre acre_40_40 (.clk(clk), .en(en), .top_left({trees[1989], lumberyards[1989]}), .top({trees[1990], lumberyards[1990]}), .top_right({trees[1991], lumberyards[1991]}), .left({trees[2039], lumberyards[2039]}), .right({trees[2041], lumberyards[2041]}), .bottom_left({trees[2089], lumberyards[2089]}), .bottom({trees[2090], lumberyards[2090]}), .bottom_right({trees[2091], lumberyards[2091]}), .init(2'b00), .state({trees[2040], lumberyards[2040]}));
acre acre_40_41 (.clk(clk), .en(en), .top_left({trees[1990], lumberyards[1990]}), .top({trees[1991], lumberyards[1991]}), .top_right({trees[1992], lumberyards[1992]}), .left({trees[2040], lumberyards[2040]}), .right({trees[2042], lumberyards[2042]}), .bottom_left({trees[2090], lumberyards[2090]}), .bottom({trees[2091], lumberyards[2091]}), .bottom_right({trees[2092], lumberyards[2092]}), .init(2'b00), .state({trees[2041], lumberyards[2041]}));
acre acre_40_42 (.clk(clk), .en(en), .top_left({trees[1991], lumberyards[1991]}), .top({trees[1992], lumberyards[1992]}), .top_right({trees[1993], lumberyards[1993]}), .left({trees[2041], lumberyards[2041]}), .right({trees[2043], lumberyards[2043]}), .bottom_left({trees[2091], lumberyards[2091]}), .bottom({trees[2092], lumberyards[2092]}), .bottom_right({trees[2093], lumberyards[2093]}), .init(2'b00), .state({trees[2042], lumberyards[2042]}));
acre acre_40_43 (.clk(clk), .en(en), .top_left({trees[1992], lumberyards[1992]}), .top({trees[1993], lumberyards[1993]}), .top_right({trees[1994], lumberyards[1994]}), .left({trees[2042], lumberyards[2042]}), .right({trees[2044], lumberyards[2044]}), .bottom_left({trees[2092], lumberyards[2092]}), .bottom({trees[2093], lumberyards[2093]}), .bottom_right({trees[2094], lumberyards[2094]}), .init(2'b01), .state({trees[2043], lumberyards[2043]}));
acre acre_40_44 (.clk(clk), .en(en), .top_left({trees[1993], lumberyards[1993]}), .top({trees[1994], lumberyards[1994]}), .top_right({trees[1995], lumberyards[1995]}), .left({trees[2043], lumberyards[2043]}), .right({trees[2045], lumberyards[2045]}), .bottom_left({trees[2093], lumberyards[2093]}), .bottom({trees[2094], lumberyards[2094]}), .bottom_right({trees[2095], lumberyards[2095]}), .init(2'b00), .state({trees[2044], lumberyards[2044]}));
acre acre_40_45 (.clk(clk), .en(en), .top_left({trees[1994], lumberyards[1994]}), .top({trees[1995], lumberyards[1995]}), .top_right({trees[1996], lumberyards[1996]}), .left({trees[2044], lumberyards[2044]}), .right({trees[2046], lumberyards[2046]}), .bottom_left({trees[2094], lumberyards[2094]}), .bottom({trees[2095], lumberyards[2095]}), .bottom_right({trees[2096], lumberyards[2096]}), .init(2'b10), .state({trees[2045], lumberyards[2045]}));
acre acre_40_46 (.clk(clk), .en(en), .top_left({trees[1995], lumberyards[1995]}), .top({trees[1996], lumberyards[1996]}), .top_right({trees[1997], lumberyards[1997]}), .left({trees[2045], lumberyards[2045]}), .right({trees[2047], lumberyards[2047]}), .bottom_left({trees[2095], lumberyards[2095]}), .bottom({trees[2096], lumberyards[2096]}), .bottom_right({trees[2097], lumberyards[2097]}), .init(2'b00), .state({trees[2046], lumberyards[2046]}));
acre acre_40_47 (.clk(clk), .en(en), .top_left({trees[1996], lumberyards[1996]}), .top({trees[1997], lumberyards[1997]}), .top_right({trees[1998], lumberyards[1998]}), .left({trees[2046], lumberyards[2046]}), .right({trees[2048], lumberyards[2048]}), .bottom_left({trees[2096], lumberyards[2096]}), .bottom({trees[2097], lumberyards[2097]}), .bottom_right({trees[2098], lumberyards[2098]}), .init(2'b00), .state({trees[2047], lumberyards[2047]}));
acre acre_40_48 (.clk(clk), .en(en), .top_left({trees[1997], lumberyards[1997]}), .top({trees[1998], lumberyards[1998]}), .top_right({trees[1999], lumberyards[1999]}), .left({trees[2047], lumberyards[2047]}), .right({trees[2049], lumberyards[2049]}), .bottom_left({trees[2097], lumberyards[2097]}), .bottom({trees[2098], lumberyards[2098]}), .bottom_right({trees[2099], lumberyards[2099]}), .init(2'b00), .state({trees[2048], lumberyards[2048]}));
acre acre_40_49 (.clk(clk), .en(en), .top_left({trees[1998], lumberyards[1998]}), .top({trees[1999], lumberyards[1999]}), .top_right(2'b0), .left({trees[2048], lumberyards[2048]}), .right(2'b0), .bottom_left({trees[2098], lumberyards[2098]}), .bottom({trees[2099], lumberyards[2099]}), .bottom_right(2'b0), .init(2'b01), .state({trees[2049], lumberyards[2049]}));
acre acre_41_0 (.clk(clk), .en(en), .top_left(2'b0), .top({trees[2000], lumberyards[2000]}), .top_right({trees[2001], lumberyards[2001]}), .left(2'b0), .right({trees[2051], lumberyards[2051]}), .bottom_left(2'b0), .bottom({trees[2100], lumberyards[2100]}), .bottom_right({trees[2101], lumberyards[2101]}), .init(2'b10), .state({trees[2050], lumberyards[2050]}));
acre acre_41_1 (.clk(clk), .en(en), .top_left({trees[2000], lumberyards[2000]}), .top({trees[2001], lumberyards[2001]}), .top_right({trees[2002], lumberyards[2002]}), .left({trees[2050], lumberyards[2050]}), .right({trees[2052], lumberyards[2052]}), .bottom_left({trees[2100], lumberyards[2100]}), .bottom({trees[2101], lumberyards[2101]}), .bottom_right({trees[2102], lumberyards[2102]}), .init(2'b00), .state({trees[2051], lumberyards[2051]}));
acre acre_41_2 (.clk(clk), .en(en), .top_left({trees[2001], lumberyards[2001]}), .top({trees[2002], lumberyards[2002]}), .top_right({trees[2003], lumberyards[2003]}), .left({trees[2051], lumberyards[2051]}), .right({trees[2053], lumberyards[2053]}), .bottom_left({trees[2101], lumberyards[2101]}), .bottom({trees[2102], lumberyards[2102]}), .bottom_right({trees[2103], lumberyards[2103]}), .init(2'b00), .state({trees[2052], lumberyards[2052]}));
acre acre_41_3 (.clk(clk), .en(en), .top_left({trees[2002], lumberyards[2002]}), .top({trees[2003], lumberyards[2003]}), .top_right({trees[2004], lumberyards[2004]}), .left({trees[2052], lumberyards[2052]}), .right({trees[2054], lumberyards[2054]}), .bottom_left({trees[2102], lumberyards[2102]}), .bottom({trees[2103], lumberyards[2103]}), .bottom_right({trees[2104], lumberyards[2104]}), .init(2'b00), .state({trees[2053], lumberyards[2053]}));
acre acre_41_4 (.clk(clk), .en(en), .top_left({trees[2003], lumberyards[2003]}), .top({trees[2004], lumberyards[2004]}), .top_right({trees[2005], lumberyards[2005]}), .left({trees[2053], lumberyards[2053]}), .right({trees[2055], lumberyards[2055]}), .bottom_left({trees[2103], lumberyards[2103]}), .bottom({trees[2104], lumberyards[2104]}), .bottom_right({trees[2105], lumberyards[2105]}), .init(2'b00), .state({trees[2054], lumberyards[2054]}));
acre acre_41_5 (.clk(clk), .en(en), .top_left({trees[2004], lumberyards[2004]}), .top({trees[2005], lumberyards[2005]}), .top_right({trees[2006], lumberyards[2006]}), .left({trees[2054], lumberyards[2054]}), .right({trees[2056], lumberyards[2056]}), .bottom_left({trees[2104], lumberyards[2104]}), .bottom({trees[2105], lumberyards[2105]}), .bottom_right({trees[2106], lumberyards[2106]}), .init(2'b00), .state({trees[2055], lumberyards[2055]}));
acre acre_41_6 (.clk(clk), .en(en), .top_left({trees[2005], lumberyards[2005]}), .top({trees[2006], lumberyards[2006]}), .top_right({trees[2007], lumberyards[2007]}), .left({trees[2055], lumberyards[2055]}), .right({trees[2057], lumberyards[2057]}), .bottom_left({trees[2105], lumberyards[2105]}), .bottom({trees[2106], lumberyards[2106]}), .bottom_right({trees[2107], lumberyards[2107]}), .init(2'b00), .state({trees[2056], lumberyards[2056]}));
acre acre_41_7 (.clk(clk), .en(en), .top_left({trees[2006], lumberyards[2006]}), .top({trees[2007], lumberyards[2007]}), .top_right({trees[2008], lumberyards[2008]}), .left({trees[2056], lumberyards[2056]}), .right({trees[2058], lumberyards[2058]}), .bottom_left({trees[2106], lumberyards[2106]}), .bottom({trees[2107], lumberyards[2107]}), .bottom_right({trees[2108], lumberyards[2108]}), .init(2'b10), .state({trees[2057], lumberyards[2057]}));
acre acre_41_8 (.clk(clk), .en(en), .top_left({trees[2007], lumberyards[2007]}), .top({trees[2008], lumberyards[2008]}), .top_right({trees[2009], lumberyards[2009]}), .left({trees[2057], lumberyards[2057]}), .right({trees[2059], lumberyards[2059]}), .bottom_left({trees[2107], lumberyards[2107]}), .bottom({trees[2108], lumberyards[2108]}), .bottom_right({trees[2109], lumberyards[2109]}), .init(2'b00), .state({trees[2058], lumberyards[2058]}));
acre acre_41_9 (.clk(clk), .en(en), .top_left({trees[2008], lumberyards[2008]}), .top({trees[2009], lumberyards[2009]}), .top_right({trees[2010], lumberyards[2010]}), .left({trees[2058], lumberyards[2058]}), .right({trees[2060], lumberyards[2060]}), .bottom_left({trees[2108], lumberyards[2108]}), .bottom({trees[2109], lumberyards[2109]}), .bottom_right({trees[2110], lumberyards[2110]}), .init(2'b00), .state({trees[2059], lumberyards[2059]}));
acre acre_41_10 (.clk(clk), .en(en), .top_left({trees[2009], lumberyards[2009]}), .top({trees[2010], lumberyards[2010]}), .top_right({trees[2011], lumberyards[2011]}), .left({trees[2059], lumberyards[2059]}), .right({trees[2061], lumberyards[2061]}), .bottom_left({trees[2109], lumberyards[2109]}), .bottom({trees[2110], lumberyards[2110]}), .bottom_right({trees[2111], lumberyards[2111]}), .init(2'b00), .state({trees[2060], lumberyards[2060]}));
acre acre_41_11 (.clk(clk), .en(en), .top_left({trees[2010], lumberyards[2010]}), .top({trees[2011], lumberyards[2011]}), .top_right({trees[2012], lumberyards[2012]}), .left({trees[2060], lumberyards[2060]}), .right({trees[2062], lumberyards[2062]}), .bottom_left({trees[2110], lumberyards[2110]}), .bottom({trees[2111], lumberyards[2111]}), .bottom_right({trees[2112], lumberyards[2112]}), .init(2'b01), .state({trees[2061], lumberyards[2061]}));
acre acre_41_12 (.clk(clk), .en(en), .top_left({trees[2011], lumberyards[2011]}), .top({trees[2012], lumberyards[2012]}), .top_right({trees[2013], lumberyards[2013]}), .left({trees[2061], lumberyards[2061]}), .right({trees[2063], lumberyards[2063]}), .bottom_left({trees[2111], lumberyards[2111]}), .bottom({trees[2112], lumberyards[2112]}), .bottom_right({trees[2113], lumberyards[2113]}), .init(2'b01), .state({trees[2062], lumberyards[2062]}));
acre acre_41_13 (.clk(clk), .en(en), .top_left({trees[2012], lumberyards[2012]}), .top({trees[2013], lumberyards[2013]}), .top_right({trees[2014], lumberyards[2014]}), .left({trees[2062], lumberyards[2062]}), .right({trees[2064], lumberyards[2064]}), .bottom_left({trees[2112], lumberyards[2112]}), .bottom({trees[2113], lumberyards[2113]}), .bottom_right({trees[2114], lumberyards[2114]}), .init(2'b01), .state({trees[2063], lumberyards[2063]}));
acre acre_41_14 (.clk(clk), .en(en), .top_left({trees[2013], lumberyards[2013]}), .top({trees[2014], lumberyards[2014]}), .top_right({trees[2015], lumberyards[2015]}), .left({trees[2063], lumberyards[2063]}), .right({trees[2065], lumberyards[2065]}), .bottom_left({trees[2113], lumberyards[2113]}), .bottom({trees[2114], lumberyards[2114]}), .bottom_right({trees[2115], lumberyards[2115]}), .init(2'b00), .state({trees[2064], lumberyards[2064]}));
acre acre_41_15 (.clk(clk), .en(en), .top_left({trees[2014], lumberyards[2014]}), .top({trees[2015], lumberyards[2015]}), .top_right({trees[2016], lumberyards[2016]}), .left({trees[2064], lumberyards[2064]}), .right({trees[2066], lumberyards[2066]}), .bottom_left({trees[2114], lumberyards[2114]}), .bottom({trees[2115], lumberyards[2115]}), .bottom_right({trees[2116], lumberyards[2116]}), .init(2'b10), .state({trees[2065], lumberyards[2065]}));
acre acre_41_16 (.clk(clk), .en(en), .top_left({trees[2015], lumberyards[2015]}), .top({trees[2016], lumberyards[2016]}), .top_right({trees[2017], lumberyards[2017]}), .left({trees[2065], lumberyards[2065]}), .right({trees[2067], lumberyards[2067]}), .bottom_left({trees[2115], lumberyards[2115]}), .bottom({trees[2116], lumberyards[2116]}), .bottom_right({trees[2117], lumberyards[2117]}), .init(2'b00), .state({trees[2066], lumberyards[2066]}));
acre acre_41_17 (.clk(clk), .en(en), .top_left({trees[2016], lumberyards[2016]}), .top({trees[2017], lumberyards[2017]}), .top_right({trees[2018], lumberyards[2018]}), .left({trees[2066], lumberyards[2066]}), .right({trees[2068], lumberyards[2068]}), .bottom_left({trees[2116], lumberyards[2116]}), .bottom({trees[2117], lumberyards[2117]}), .bottom_right({trees[2118], lumberyards[2118]}), .init(2'b00), .state({trees[2067], lumberyards[2067]}));
acre acre_41_18 (.clk(clk), .en(en), .top_left({trees[2017], lumberyards[2017]}), .top({trees[2018], lumberyards[2018]}), .top_right({trees[2019], lumberyards[2019]}), .left({trees[2067], lumberyards[2067]}), .right({trees[2069], lumberyards[2069]}), .bottom_left({trees[2117], lumberyards[2117]}), .bottom({trees[2118], lumberyards[2118]}), .bottom_right({trees[2119], lumberyards[2119]}), .init(2'b01), .state({trees[2068], lumberyards[2068]}));
acre acre_41_19 (.clk(clk), .en(en), .top_left({trees[2018], lumberyards[2018]}), .top({trees[2019], lumberyards[2019]}), .top_right({trees[2020], lumberyards[2020]}), .left({trees[2068], lumberyards[2068]}), .right({trees[2070], lumberyards[2070]}), .bottom_left({trees[2118], lumberyards[2118]}), .bottom({trees[2119], lumberyards[2119]}), .bottom_right({trees[2120], lumberyards[2120]}), .init(2'b00), .state({trees[2069], lumberyards[2069]}));
acre acre_41_20 (.clk(clk), .en(en), .top_left({trees[2019], lumberyards[2019]}), .top({trees[2020], lumberyards[2020]}), .top_right({trees[2021], lumberyards[2021]}), .left({trees[2069], lumberyards[2069]}), .right({trees[2071], lumberyards[2071]}), .bottom_left({trees[2119], lumberyards[2119]}), .bottom({trees[2120], lumberyards[2120]}), .bottom_right({trees[2121], lumberyards[2121]}), .init(2'b10), .state({trees[2070], lumberyards[2070]}));
acre acre_41_21 (.clk(clk), .en(en), .top_left({trees[2020], lumberyards[2020]}), .top({trees[2021], lumberyards[2021]}), .top_right({trees[2022], lumberyards[2022]}), .left({trees[2070], lumberyards[2070]}), .right({trees[2072], lumberyards[2072]}), .bottom_left({trees[2120], lumberyards[2120]}), .bottom({trees[2121], lumberyards[2121]}), .bottom_right({trees[2122], lumberyards[2122]}), .init(2'b01), .state({trees[2071], lumberyards[2071]}));
acre acre_41_22 (.clk(clk), .en(en), .top_left({trees[2021], lumberyards[2021]}), .top({trees[2022], lumberyards[2022]}), .top_right({trees[2023], lumberyards[2023]}), .left({trees[2071], lumberyards[2071]}), .right({trees[2073], lumberyards[2073]}), .bottom_left({trees[2121], lumberyards[2121]}), .bottom({trees[2122], lumberyards[2122]}), .bottom_right({trees[2123], lumberyards[2123]}), .init(2'b01), .state({trees[2072], lumberyards[2072]}));
acre acre_41_23 (.clk(clk), .en(en), .top_left({trees[2022], lumberyards[2022]}), .top({trees[2023], lumberyards[2023]}), .top_right({trees[2024], lumberyards[2024]}), .left({trees[2072], lumberyards[2072]}), .right({trees[2074], lumberyards[2074]}), .bottom_left({trees[2122], lumberyards[2122]}), .bottom({trees[2123], lumberyards[2123]}), .bottom_right({trees[2124], lumberyards[2124]}), .init(2'b00), .state({trees[2073], lumberyards[2073]}));
acre acre_41_24 (.clk(clk), .en(en), .top_left({trees[2023], lumberyards[2023]}), .top({trees[2024], lumberyards[2024]}), .top_right({trees[2025], lumberyards[2025]}), .left({trees[2073], lumberyards[2073]}), .right({trees[2075], lumberyards[2075]}), .bottom_left({trees[2123], lumberyards[2123]}), .bottom({trees[2124], lumberyards[2124]}), .bottom_right({trees[2125], lumberyards[2125]}), .init(2'b00), .state({trees[2074], lumberyards[2074]}));
acre acre_41_25 (.clk(clk), .en(en), .top_left({trees[2024], lumberyards[2024]}), .top({trees[2025], lumberyards[2025]}), .top_right({trees[2026], lumberyards[2026]}), .left({trees[2074], lumberyards[2074]}), .right({trees[2076], lumberyards[2076]}), .bottom_left({trees[2124], lumberyards[2124]}), .bottom({trees[2125], lumberyards[2125]}), .bottom_right({trees[2126], lumberyards[2126]}), .init(2'b10), .state({trees[2075], lumberyards[2075]}));
acre acre_41_26 (.clk(clk), .en(en), .top_left({trees[2025], lumberyards[2025]}), .top({trees[2026], lumberyards[2026]}), .top_right({trees[2027], lumberyards[2027]}), .left({trees[2075], lumberyards[2075]}), .right({trees[2077], lumberyards[2077]}), .bottom_left({trees[2125], lumberyards[2125]}), .bottom({trees[2126], lumberyards[2126]}), .bottom_right({trees[2127], lumberyards[2127]}), .init(2'b00), .state({trees[2076], lumberyards[2076]}));
acre acre_41_27 (.clk(clk), .en(en), .top_left({trees[2026], lumberyards[2026]}), .top({trees[2027], lumberyards[2027]}), .top_right({trees[2028], lumberyards[2028]}), .left({trees[2076], lumberyards[2076]}), .right({trees[2078], lumberyards[2078]}), .bottom_left({trees[2126], lumberyards[2126]}), .bottom({trees[2127], lumberyards[2127]}), .bottom_right({trees[2128], lumberyards[2128]}), .init(2'b00), .state({trees[2077], lumberyards[2077]}));
acre acre_41_28 (.clk(clk), .en(en), .top_left({trees[2027], lumberyards[2027]}), .top({trees[2028], lumberyards[2028]}), .top_right({trees[2029], lumberyards[2029]}), .left({trees[2077], lumberyards[2077]}), .right({trees[2079], lumberyards[2079]}), .bottom_left({trees[2127], lumberyards[2127]}), .bottom({trees[2128], lumberyards[2128]}), .bottom_right({trees[2129], lumberyards[2129]}), .init(2'b00), .state({trees[2078], lumberyards[2078]}));
acre acre_41_29 (.clk(clk), .en(en), .top_left({trees[2028], lumberyards[2028]}), .top({trees[2029], lumberyards[2029]}), .top_right({trees[2030], lumberyards[2030]}), .left({trees[2078], lumberyards[2078]}), .right({trees[2080], lumberyards[2080]}), .bottom_left({trees[2128], lumberyards[2128]}), .bottom({trees[2129], lumberyards[2129]}), .bottom_right({trees[2130], lumberyards[2130]}), .init(2'b00), .state({trees[2079], lumberyards[2079]}));
acre acre_41_30 (.clk(clk), .en(en), .top_left({trees[2029], lumberyards[2029]}), .top({trees[2030], lumberyards[2030]}), .top_right({trees[2031], lumberyards[2031]}), .left({trees[2079], lumberyards[2079]}), .right({trees[2081], lumberyards[2081]}), .bottom_left({trees[2129], lumberyards[2129]}), .bottom({trees[2130], lumberyards[2130]}), .bottom_right({trees[2131], lumberyards[2131]}), .init(2'b00), .state({trees[2080], lumberyards[2080]}));
acre acre_41_31 (.clk(clk), .en(en), .top_left({trees[2030], lumberyards[2030]}), .top({trees[2031], lumberyards[2031]}), .top_right({trees[2032], lumberyards[2032]}), .left({trees[2080], lumberyards[2080]}), .right({trees[2082], lumberyards[2082]}), .bottom_left({trees[2130], lumberyards[2130]}), .bottom({trees[2131], lumberyards[2131]}), .bottom_right({trees[2132], lumberyards[2132]}), .init(2'b00), .state({trees[2081], lumberyards[2081]}));
acre acre_41_32 (.clk(clk), .en(en), .top_left({trees[2031], lumberyards[2031]}), .top({trees[2032], lumberyards[2032]}), .top_right({trees[2033], lumberyards[2033]}), .left({trees[2081], lumberyards[2081]}), .right({trees[2083], lumberyards[2083]}), .bottom_left({trees[2131], lumberyards[2131]}), .bottom({trees[2132], lumberyards[2132]}), .bottom_right({trees[2133], lumberyards[2133]}), .init(2'b00), .state({trees[2082], lumberyards[2082]}));
acre acre_41_33 (.clk(clk), .en(en), .top_left({trees[2032], lumberyards[2032]}), .top({trees[2033], lumberyards[2033]}), .top_right({trees[2034], lumberyards[2034]}), .left({trees[2082], lumberyards[2082]}), .right({trees[2084], lumberyards[2084]}), .bottom_left({trees[2132], lumberyards[2132]}), .bottom({trees[2133], lumberyards[2133]}), .bottom_right({trees[2134], lumberyards[2134]}), .init(2'b10), .state({trees[2083], lumberyards[2083]}));
acre acre_41_34 (.clk(clk), .en(en), .top_left({trees[2033], lumberyards[2033]}), .top({trees[2034], lumberyards[2034]}), .top_right({trees[2035], lumberyards[2035]}), .left({trees[2083], lumberyards[2083]}), .right({trees[2085], lumberyards[2085]}), .bottom_left({trees[2133], lumberyards[2133]}), .bottom({trees[2134], lumberyards[2134]}), .bottom_right({trees[2135], lumberyards[2135]}), .init(2'b00), .state({trees[2084], lumberyards[2084]}));
acre acre_41_35 (.clk(clk), .en(en), .top_left({trees[2034], lumberyards[2034]}), .top({trees[2035], lumberyards[2035]}), .top_right({trees[2036], lumberyards[2036]}), .left({trees[2084], lumberyards[2084]}), .right({trees[2086], lumberyards[2086]}), .bottom_left({trees[2134], lumberyards[2134]}), .bottom({trees[2135], lumberyards[2135]}), .bottom_right({trees[2136], lumberyards[2136]}), .init(2'b10), .state({trees[2085], lumberyards[2085]}));
acre acre_41_36 (.clk(clk), .en(en), .top_left({trees[2035], lumberyards[2035]}), .top({trees[2036], lumberyards[2036]}), .top_right({trees[2037], lumberyards[2037]}), .left({trees[2085], lumberyards[2085]}), .right({trees[2087], lumberyards[2087]}), .bottom_left({trees[2135], lumberyards[2135]}), .bottom({trees[2136], lumberyards[2136]}), .bottom_right({trees[2137], lumberyards[2137]}), .init(2'b00), .state({trees[2086], lumberyards[2086]}));
acre acre_41_37 (.clk(clk), .en(en), .top_left({trees[2036], lumberyards[2036]}), .top({trees[2037], lumberyards[2037]}), .top_right({trees[2038], lumberyards[2038]}), .left({trees[2086], lumberyards[2086]}), .right({trees[2088], lumberyards[2088]}), .bottom_left({trees[2136], lumberyards[2136]}), .bottom({trees[2137], lumberyards[2137]}), .bottom_right({trees[2138], lumberyards[2138]}), .init(2'b01), .state({trees[2087], lumberyards[2087]}));
acre acre_41_38 (.clk(clk), .en(en), .top_left({trees[2037], lumberyards[2037]}), .top({trees[2038], lumberyards[2038]}), .top_right({trees[2039], lumberyards[2039]}), .left({trees[2087], lumberyards[2087]}), .right({trees[2089], lumberyards[2089]}), .bottom_left({trees[2137], lumberyards[2137]}), .bottom({trees[2138], lumberyards[2138]}), .bottom_right({trees[2139], lumberyards[2139]}), .init(2'b00), .state({trees[2088], lumberyards[2088]}));
acre acre_41_39 (.clk(clk), .en(en), .top_left({trees[2038], lumberyards[2038]}), .top({trees[2039], lumberyards[2039]}), .top_right({trees[2040], lumberyards[2040]}), .left({trees[2088], lumberyards[2088]}), .right({trees[2090], lumberyards[2090]}), .bottom_left({trees[2138], lumberyards[2138]}), .bottom({trees[2139], lumberyards[2139]}), .bottom_right({trees[2140], lumberyards[2140]}), .init(2'b00), .state({trees[2089], lumberyards[2089]}));
acre acre_41_40 (.clk(clk), .en(en), .top_left({trees[2039], lumberyards[2039]}), .top({trees[2040], lumberyards[2040]}), .top_right({trees[2041], lumberyards[2041]}), .left({trees[2089], lumberyards[2089]}), .right({trees[2091], lumberyards[2091]}), .bottom_left({trees[2139], lumberyards[2139]}), .bottom({trees[2140], lumberyards[2140]}), .bottom_right({trees[2141], lumberyards[2141]}), .init(2'b00), .state({trees[2090], lumberyards[2090]}));
acre acre_41_41 (.clk(clk), .en(en), .top_left({trees[2040], lumberyards[2040]}), .top({trees[2041], lumberyards[2041]}), .top_right({trees[2042], lumberyards[2042]}), .left({trees[2090], lumberyards[2090]}), .right({trees[2092], lumberyards[2092]}), .bottom_left({trees[2140], lumberyards[2140]}), .bottom({trees[2141], lumberyards[2141]}), .bottom_right({trees[2142], lumberyards[2142]}), .init(2'b10), .state({trees[2091], lumberyards[2091]}));
acre acre_41_42 (.clk(clk), .en(en), .top_left({trees[2041], lumberyards[2041]}), .top({trees[2042], lumberyards[2042]}), .top_right({trees[2043], lumberyards[2043]}), .left({trees[2091], lumberyards[2091]}), .right({trees[2093], lumberyards[2093]}), .bottom_left({trees[2141], lumberyards[2141]}), .bottom({trees[2142], lumberyards[2142]}), .bottom_right({trees[2143], lumberyards[2143]}), .init(2'b00), .state({trees[2092], lumberyards[2092]}));
acre acre_41_43 (.clk(clk), .en(en), .top_left({trees[2042], lumberyards[2042]}), .top({trees[2043], lumberyards[2043]}), .top_right({trees[2044], lumberyards[2044]}), .left({trees[2092], lumberyards[2092]}), .right({trees[2094], lumberyards[2094]}), .bottom_left({trees[2142], lumberyards[2142]}), .bottom({trees[2143], lumberyards[2143]}), .bottom_right({trees[2144], lumberyards[2144]}), .init(2'b00), .state({trees[2093], lumberyards[2093]}));
acre acre_41_44 (.clk(clk), .en(en), .top_left({trees[2043], lumberyards[2043]}), .top({trees[2044], lumberyards[2044]}), .top_right({trees[2045], lumberyards[2045]}), .left({trees[2093], lumberyards[2093]}), .right({trees[2095], lumberyards[2095]}), .bottom_left({trees[2143], lumberyards[2143]}), .bottom({trees[2144], lumberyards[2144]}), .bottom_right({trees[2145], lumberyards[2145]}), .init(2'b10), .state({trees[2094], lumberyards[2094]}));
acre acre_41_45 (.clk(clk), .en(en), .top_left({trees[2044], lumberyards[2044]}), .top({trees[2045], lumberyards[2045]}), .top_right({trees[2046], lumberyards[2046]}), .left({trees[2094], lumberyards[2094]}), .right({trees[2096], lumberyards[2096]}), .bottom_left({trees[2144], lumberyards[2144]}), .bottom({trees[2145], lumberyards[2145]}), .bottom_right({trees[2146], lumberyards[2146]}), .init(2'b00), .state({trees[2095], lumberyards[2095]}));
acre acre_41_46 (.clk(clk), .en(en), .top_left({trees[2045], lumberyards[2045]}), .top({trees[2046], lumberyards[2046]}), .top_right({trees[2047], lumberyards[2047]}), .left({trees[2095], lumberyards[2095]}), .right({trees[2097], lumberyards[2097]}), .bottom_left({trees[2145], lumberyards[2145]}), .bottom({trees[2146], lumberyards[2146]}), .bottom_right({trees[2147], lumberyards[2147]}), .init(2'b01), .state({trees[2096], lumberyards[2096]}));
acre acre_41_47 (.clk(clk), .en(en), .top_left({trees[2046], lumberyards[2046]}), .top({trees[2047], lumberyards[2047]}), .top_right({trees[2048], lumberyards[2048]}), .left({trees[2096], lumberyards[2096]}), .right({trees[2098], lumberyards[2098]}), .bottom_left({trees[2146], lumberyards[2146]}), .bottom({trees[2147], lumberyards[2147]}), .bottom_right({trees[2148], lumberyards[2148]}), .init(2'b00), .state({trees[2097], lumberyards[2097]}));
acre acre_41_48 (.clk(clk), .en(en), .top_left({trees[2047], lumberyards[2047]}), .top({trees[2048], lumberyards[2048]}), .top_right({trees[2049], lumberyards[2049]}), .left({trees[2097], lumberyards[2097]}), .right({trees[2099], lumberyards[2099]}), .bottom_left({trees[2147], lumberyards[2147]}), .bottom({trees[2148], lumberyards[2148]}), .bottom_right({trees[2149], lumberyards[2149]}), .init(2'b01), .state({trees[2098], lumberyards[2098]}));
acre acre_41_49 (.clk(clk), .en(en), .top_left({trees[2048], lumberyards[2048]}), .top({trees[2049], lumberyards[2049]}), .top_right(2'b0), .left({trees[2098], lumberyards[2098]}), .right(2'b0), .bottom_left({trees[2148], lumberyards[2148]}), .bottom({trees[2149], lumberyards[2149]}), .bottom_right(2'b0), .init(2'b01), .state({trees[2099], lumberyards[2099]}));
acre acre_42_0 (.clk(clk), .en(en), .top_left(2'b0), .top({trees[2050], lumberyards[2050]}), .top_right({trees[2051], lumberyards[2051]}), .left(2'b0), .right({trees[2101], lumberyards[2101]}), .bottom_left(2'b0), .bottom({trees[2150], lumberyards[2150]}), .bottom_right({trees[2151], lumberyards[2151]}), .init(2'b10), .state({trees[2100], lumberyards[2100]}));
acre acre_42_1 (.clk(clk), .en(en), .top_left({trees[2050], lumberyards[2050]}), .top({trees[2051], lumberyards[2051]}), .top_right({trees[2052], lumberyards[2052]}), .left({trees[2100], lumberyards[2100]}), .right({trees[2102], lumberyards[2102]}), .bottom_left({trees[2150], lumberyards[2150]}), .bottom({trees[2151], lumberyards[2151]}), .bottom_right({trees[2152], lumberyards[2152]}), .init(2'b00), .state({trees[2101], lumberyards[2101]}));
acre acre_42_2 (.clk(clk), .en(en), .top_left({trees[2051], lumberyards[2051]}), .top({trees[2052], lumberyards[2052]}), .top_right({trees[2053], lumberyards[2053]}), .left({trees[2101], lumberyards[2101]}), .right({trees[2103], lumberyards[2103]}), .bottom_left({trees[2151], lumberyards[2151]}), .bottom({trees[2152], lumberyards[2152]}), .bottom_right({trees[2153], lumberyards[2153]}), .init(2'b00), .state({trees[2102], lumberyards[2102]}));
acre acre_42_3 (.clk(clk), .en(en), .top_left({trees[2052], lumberyards[2052]}), .top({trees[2053], lumberyards[2053]}), .top_right({trees[2054], lumberyards[2054]}), .left({trees[2102], lumberyards[2102]}), .right({trees[2104], lumberyards[2104]}), .bottom_left({trees[2152], lumberyards[2152]}), .bottom({trees[2153], lumberyards[2153]}), .bottom_right({trees[2154], lumberyards[2154]}), .init(2'b00), .state({trees[2103], lumberyards[2103]}));
acre acre_42_4 (.clk(clk), .en(en), .top_left({trees[2053], lumberyards[2053]}), .top({trees[2054], lumberyards[2054]}), .top_right({trees[2055], lumberyards[2055]}), .left({trees[2103], lumberyards[2103]}), .right({trees[2105], lumberyards[2105]}), .bottom_left({trees[2153], lumberyards[2153]}), .bottom({trees[2154], lumberyards[2154]}), .bottom_right({trees[2155], lumberyards[2155]}), .init(2'b00), .state({trees[2104], lumberyards[2104]}));
acre acre_42_5 (.clk(clk), .en(en), .top_left({trees[2054], lumberyards[2054]}), .top({trees[2055], lumberyards[2055]}), .top_right({trees[2056], lumberyards[2056]}), .left({trees[2104], lumberyards[2104]}), .right({trees[2106], lumberyards[2106]}), .bottom_left({trees[2154], lumberyards[2154]}), .bottom({trees[2155], lumberyards[2155]}), .bottom_right({trees[2156], lumberyards[2156]}), .init(2'b00), .state({trees[2105], lumberyards[2105]}));
acre acre_42_6 (.clk(clk), .en(en), .top_left({trees[2055], lumberyards[2055]}), .top({trees[2056], lumberyards[2056]}), .top_right({trees[2057], lumberyards[2057]}), .left({trees[2105], lumberyards[2105]}), .right({trees[2107], lumberyards[2107]}), .bottom_left({trees[2155], lumberyards[2155]}), .bottom({trees[2156], lumberyards[2156]}), .bottom_right({trees[2157], lumberyards[2157]}), .init(2'b00), .state({trees[2106], lumberyards[2106]}));
acre acre_42_7 (.clk(clk), .en(en), .top_left({trees[2056], lumberyards[2056]}), .top({trees[2057], lumberyards[2057]}), .top_right({trees[2058], lumberyards[2058]}), .left({trees[2106], lumberyards[2106]}), .right({trees[2108], lumberyards[2108]}), .bottom_left({trees[2156], lumberyards[2156]}), .bottom({trees[2157], lumberyards[2157]}), .bottom_right({trees[2158], lumberyards[2158]}), .init(2'b01), .state({trees[2107], lumberyards[2107]}));
acre acre_42_8 (.clk(clk), .en(en), .top_left({trees[2057], lumberyards[2057]}), .top({trees[2058], lumberyards[2058]}), .top_right({trees[2059], lumberyards[2059]}), .left({trees[2107], lumberyards[2107]}), .right({trees[2109], lumberyards[2109]}), .bottom_left({trees[2157], lumberyards[2157]}), .bottom({trees[2158], lumberyards[2158]}), .bottom_right({trees[2159], lumberyards[2159]}), .init(2'b00), .state({trees[2108], lumberyards[2108]}));
acre acre_42_9 (.clk(clk), .en(en), .top_left({trees[2058], lumberyards[2058]}), .top({trees[2059], lumberyards[2059]}), .top_right({trees[2060], lumberyards[2060]}), .left({trees[2108], lumberyards[2108]}), .right({trees[2110], lumberyards[2110]}), .bottom_left({trees[2158], lumberyards[2158]}), .bottom({trees[2159], lumberyards[2159]}), .bottom_right({trees[2160], lumberyards[2160]}), .init(2'b00), .state({trees[2109], lumberyards[2109]}));
acre acre_42_10 (.clk(clk), .en(en), .top_left({trees[2059], lumberyards[2059]}), .top({trees[2060], lumberyards[2060]}), .top_right({trees[2061], lumberyards[2061]}), .left({trees[2109], lumberyards[2109]}), .right({trees[2111], lumberyards[2111]}), .bottom_left({trees[2159], lumberyards[2159]}), .bottom({trees[2160], lumberyards[2160]}), .bottom_right({trees[2161], lumberyards[2161]}), .init(2'b00), .state({trees[2110], lumberyards[2110]}));
acre acre_42_11 (.clk(clk), .en(en), .top_left({trees[2060], lumberyards[2060]}), .top({trees[2061], lumberyards[2061]}), .top_right({trees[2062], lumberyards[2062]}), .left({trees[2110], lumberyards[2110]}), .right({trees[2112], lumberyards[2112]}), .bottom_left({trees[2160], lumberyards[2160]}), .bottom({trees[2161], lumberyards[2161]}), .bottom_right({trees[2162], lumberyards[2162]}), .init(2'b00), .state({trees[2111], lumberyards[2111]}));
acre acre_42_12 (.clk(clk), .en(en), .top_left({trees[2061], lumberyards[2061]}), .top({trees[2062], lumberyards[2062]}), .top_right({trees[2063], lumberyards[2063]}), .left({trees[2111], lumberyards[2111]}), .right({trees[2113], lumberyards[2113]}), .bottom_left({trees[2161], lumberyards[2161]}), .bottom({trees[2162], lumberyards[2162]}), .bottom_right({trees[2163], lumberyards[2163]}), .init(2'b00), .state({trees[2112], lumberyards[2112]}));
acre acre_42_13 (.clk(clk), .en(en), .top_left({trees[2062], lumberyards[2062]}), .top({trees[2063], lumberyards[2063]}), .top_right({trees[2064], lumberyards[2064]}), .left({trees[2112], lumberyards[2112]}), .right({trees[2114], lumberyards[2114]}), .bottom_left({trees[2162], lumberyards[2162]}), .bottom({trees[2163], lumberyards[2163]}), .bottom_right({trees[2164], lumberyards[2164]}), .init(2'b01), .state({trees[2113], lumberyards[2113]}));
acre acre_42_14 (.clk(clk), .en(en), .top_left({trees[2063], lumberyards[2063]}), .top({trees[2064], lumberyards[2064]}), .top_right({trees[2065], lumberyards[2065]}), .left({trees[2113], lumberyards[2113]}), .right({trees[2115], lumberyards[2115]}), .bottom_left({trees[2163], lumberyards[2163]}), .bottom({trees[2164], lumberyards[2164]}), .bottom_right({trees[2165], lumberyards[2165]}), .init(2'b00), .state({trees[2114], lumberyards[2114]}));
acre acre_42_15 (.clk(clk), .en(en), .top_left({trees[2064], lumberyards[2064]}), .top({trees[2065], lumberyards[2065]}), .top_right({trees[2066], lumberyards[2066]}), .left({trees[2114], lumberyards[2114]}), .right({trees[2116], lumberyards[2116]}), .bottom_left({trees[2164], lumberyards[2164]}), .bottom({trees[2165], lumberyards[2165]}), .bottom_right({trees[2166], lumberyards[2166]}), .init(2'b00), .state({trees[2115], lumberyards[2115]}));
acre acre_42_16 (.clk(clk), .en(en), .top_left({trees[2065], lumberyards[2065]}), .top({trees[2066], lumberyards[2066]}), .top_right({trees[2067], lumberyards[2067]}), .left({trees[2115], lumberyards[2115]}), .right({trees[2117], lumberyards[2117]}), .bottom_left({trees[2165], lumberyards[2165]}), .bottom({trees[2166], lumberyards[2166]}), .bottom_right({trees[2167], lumberyards[2167]}), .init(2'b01), .state({trees[2116], lumberyards[2116]}));
acre acre_42_17 (.clk(clk), .en(en), .top_left({trees[2066], lumberyards[2066]}), .top({trees[2067], lumberyards[2067]}), .top_right({trees[2068], lumberyards[2068]}), .left({trees[2116], lumberyards[2116]}), .right({trees[2118], lumberyards[2118]}), .bottom_left({trees[2166], lumberyards[2166]}), .bottom({trees[2167], lumberyards[2167]}), .bottom_right({trees[2168], lumberyards[2168]}), .init(2'b10), .state({trees[2117], lumberyards[2117]}));
acre acre_42_18 (.clk(clk), .en(en), .top_left({trees[2067], lumberyards[2067]}), .top({trees[2068], lumberyards[2068]}), .top_right({trees[2069], lumberyards[2069]}), .left({trees[2117], lumberyards[2117]}), .right({trees[2119], lumberyards[2119]}), .bottom_left({trees[2167], lumberyards[2167]}), .bottom({trees[2168], lumberyards[2168]}), .bottom_right({trees[2169], lumberyards[2169]}), .init(2'b10), .state({trees[2118], lumberyards[2118]}));
acre acre_42_19 (.clk(clk), .en(en), .top_left({trees[2068], lumberyards[2068]}), .top({trees[2069], lumberyards[2069]}), .top_right({trees[2070], lumberyards[2070]}), .left({trees[2118], lumberyards[2118]}), .right({trees[2120], lumberyards[2120]}), .bottom_left({trees[2168], lumberyards[2168]}), .bottom({trees[2169], lumberyards[2169]}), .bottom_right({trees[2170], lumberyards[2170]}), .init(2'b00), .state({trees[2119], lumberyards[2119]}));
acre acre_42_20 (.clk(clk), .en(en), .top_left({trees[2069], lumberyards[2069]}), .top({trees[2070], lumberyards[2070]}), .top_right({trees[2071], lumberyards[2071]}), .left({trees[2119], lumberyards[2119]}), .right({trees[2121], lumberyards[2121]}), .bottom_left({trees[2169], lumberyards[2169]}), .bottom({trees[2170], lumberyards[2170]}), .bottom_right({trees[2171], lumberyards[2171]}), .init(2'b00), .state({trees[2120], lumberyards[2120]}));
acre acre_42_21 (.clk(clk), .en(en), .top_left({trees[2070], lumberyards[2070]}), .top({trees[2071], lumberyards[2071]}), .top_right({trees[2072], lumberyards[2072]}), .left({trees[2120], lumberyards[2120]}), .right({trees[2122], lumberyards[2122]}), .bottom_left({trees[2170], lumberyards[2170]}), .bottom({trees[2171], lumberyards[2171]}), .bottom_right({trees[2172], lumberyards[2172]}), .init(2'b00), .state({trees[2121], lumberyards[2121]}));
acre acre_42_22 (.clk(clk), .en(en), .top_left({trees[2071], lumberyards[2071]}), .top({trees[2072], lumberyards[2072]}), .top_right({trees[2073], lumberyards[2073]}), .left({trees[2121], lumberyards[2121]}), .right({trees[2123], lumberyards[2123]}), .bottom_left({trees[2171], lumberyards[2171]}), .bottom({trees[2172], lumberyards[2172]}), .bottom_right({trees[2173], lumberyards[2173]}), .init(2'b01), .state({trees[2122], lumberyards[2122]}));
acre acre_42_23 (.clk(clk), .en(en), .top_left({trees[2072], lumberyards[2072]}), .top({trees[2073], lumberyards[2073]}), .top_right({trees[2074], lumberyards[2074]}), .left({trees[2122], lumberyards[2122]}), .right({trees[2124], lumberyards[2124]}), .bottom_left({trees[2172], lumberyards[2172]}), .bottom({trees[2173], lumberyards[2173]}), .bottom_right({trees[2174], lumberyards[2174]}), .init(2'b01), .state({trees[2123], lumberyards[2123]}));
acre acre_42_24 (.clk(clk), .en(en), .top_left({trees[2073], lumberyards[2073]}), .top({trees[2074], lumberyards[2074]}), .top_right({trees[2075], lumberyards[2075]}), .left({trees[2123], lumberyards[2123]}), .right({trees[2125], lumberyards[2125]}), .bottom_left({trees[2173], lumberyards[2173]}), .bottom({trees[2174], lumberyards[2174]}), .bottom_right({trees[2175], lumberyards[2175]}), .init(2'b01), .state({trees[2124], lumberyards[2124]}));
acre acre_42_25 (.clk(clk), .en(en), .top_left({trees[2074], lumberyards[2074]}), .top({trees[2075], lumberyards[2075]}), .top_right({trees[2076], lumberyards[2076]}), .left({trees[2124], lumberyards[2124]}), .right({trees[2126], lumberyards[2126]}), .bottom_left({trees[2174], lumberyards[2174]}), .bottom({trees[2175], lumberyards[2175]}), .bottom_right({trees[2176], lumberyards[2176]}), .init(2'b00), .state({trees[2125], lumberyards[2125]}));
acre acre_42_26 (.clk(clk), .en(en), .top_left({trees[2075], lumberyards[2075]}), .top({trees[2076], lumberyards[2076]}), .top_right({trees[2077], lumberyards[2077]}), .left({trees[2125], lumberyards[2125]}), .right({trees[2127], lumberyards[2127]}), .bottom_left({trees[2175], lumberyards[2175]}), .bottom({trees[2176], lumberyards[2176]}), .bottom_right({trees[2177], lumberyards[2177]}), .init(2'b00), .state({trees[2126], lumberyards[2126]}));
acre acre_42_27 (.clk(clk), .en(en), .top_left({trees[2076], lumberyards[2076]}), .top({trees[2077], lumberyards[2077]}), .top_right({trees[2078], lumberyards[2078]}), .left({trees[2126], lumberyards[2126]}), .right({trees[2128], lumberyards[2128]}), .bottom_left({trees[2176], lumberyards[2176]}), .bottom({trees[2177], lumberyards[2177]}), .bottom_right({trees[2178], lumberyards[2178]}), .init(2'b01), .state({trees[2127], lumberyards[2127]}));
acre acre_42_28 (.clk(clk), .en(en), .top_left({trees[2077], lumberyards[2077]}), .top({trees[2078], lumberyards[2078]}), .top_right({trees[2079], lumberyards[2079]}), .left({trees[2127], lumberyards[2127]}), .right({trees[2129], lumberyards[2129]}), .bottom_left({trees[2177], lumberyards[2177]}), .bottom({trees[2178], lumberyards[2178]}), .bottom_right({trees[2179], lumberyards[2179]}), .init(2'b00), .state({trees[2128], lumberyards[2128]}));
acre acre_42_29 (.clk(clk), .en(en), .top_left({trees[2078], lumberyards[2078]}), .top({trees[2079], lumberyards[2079]}), .top_right({trees[2080], lumberyards[2080]}), .left({trees[2128], lumberyards[2128]}), .right({trees[2130], lumberyards[2130]}), .bottom_left({trees[2178], lumberyards[2178]}), .bottom({trees[2179], lumberyards[2179]}), .bottom_right({trees[2180], lumberyards[2180]}), .init(2'b00), .state({trees[2129], lumberyards[2129]}));
acre acre_42_30 (.clk(clk), .en(en), .top_left({trees[2079], lumberyards[2079]}), .top({trees[2080], lumberyards[2080]}), .top_right({trees[2081], lumberyards[2081]}), .left({trees[2129], lumberyards[2129]}), .right({trees[2131], lumberyards[2131]}), .bottom_left({trees[2179], lumberyards[2179]}), .bottom({trees[2180], lumberyards[2180]}), .bottom_right({trees[2181], lumberyards[2181]}), .init(2'b10), .state({trees[2130], lumberyards[2130]}));
acre acre_42_31 (.clk(clk), .en(en), .top_left({trees[2080], lumberyards[2080]}), .top({trees[2081], lumberyards[2081]}), .top_right({trees[2082], lumberyards[2082]}), .left({trees[2130], lumberyards[2130]}), .right({trees[2132], lumberyards[2132]}), .bottom_left({trees[2180], lumberyards[2180]}), .bottom({trees[2181], lumberyards[2181]}), .bottom_right({trees[2182], lumberyards[2182]}), .init(2'b00), .state({trees[2131], lumberyards[2131]}));
acre acre_42_32 (.clk(clk), .en(en), .top_left({trees[2081], lumberyards[2081]}), .top({trees[2082], lumberyards[2082]}), .top_right({trees[2083], lumberyards[2083]}), .left({trees[2131], lumberyards[2131]}), .right({trees[2133], lumberyards[2133]}), .bottom_left({trees[2181], lumberyards[2181]}), .bottom({trees[2182], lumberyards[2182]}), .bottom_right({trees[2183], lumberyards[2183]}), .init(2'b10), .state({trees[2132], lumberyards[2132]}));
acre acre_42_33 (.clk(clk), .en(en), .top_left({trees[2082], lumberyards[2082]}), .top({trees[2083], lumberyards[2083]}), .top_right({trees[2084], lumberyards[2084]}), .left({trees[2132], lumberyards[2132]}), .right({trees[2134], lumberyards[2134]}), .bottom_left({trees[2182], lumberyards[2182]}), .bottom({trees[2183], lumberyards[2183]}), .bottom_right({trees[2184], lumberyards[2184]}), .init(2'b00), .state({trees[2133], lumberyards[2133]}));
acre acre_42_34 (.clk(clk), .en(en), .top_left({trees[2083], lumberyards[2083]}), .top({trees[2084], lumberyards[2084]}), .top_right({trees[2085], lumberyards[2085]}), .left({trees[2133], lumberyards[2133]}), .right({trees[2135], lumberyards[2135]}), .bottom_left({trees[2183], lumberyards[2183]}), .bottom({trees[2184], lumberyards[2184]}), .bottom_right({trees[2185], lumberyards[2185]}), .init(2'b00), .state({trees[2134], lumberyards[2134]}));
acre acre_42_35 (.clk(clk), .en(en), .top_left({trees[2084], lumberyards[2084]}), .top({trees[2085], lumberyards[2085]}), .top_right({trees[2086], lumberyards[2086]}), .left({trees[2134], lumberyards[2134]}), .right({trees[2136], lumberyards[2136]}), .bottom_left({trees[2184], lumberyards[2184]}), .bottom({trees[2185], lumberyards[2185]}), .bottom_right({trees[2186], lumberyards[2186]}), .init(2'b01), .state({trees[2135], lumberyards[2135]}));
acre acre_42_36 (.clk(clk), .en(en), .top_left({trees[2085], lumberyards[2085]}), .top({trees[2086], lumberyards[2086]}), .top_right({trees[2087], lumberyards[2087]}), .left({trees[2135], lumberyards[2135]}), .right({trees[2137], lumberyards[2137]}), .bottom_left({trees[2185], lumberyards[2185]}), .bottom({trees[2186], lumberyards[2186]}), .bottom_right({trees[2187], lumberyards[2187]}), .init(2'b00), .state({trees[2136], lumberyards[2136]}));
acre acre_42_37 (.clk(clk), .en(en), .top_left({trees[2086], lumberyards[2086]}), .top({trees[2087], lumberyards[2087]}), .top_right({trees[2088], lumberyards[2088]}), .left({trees[2136], lumberyards[2136]}), .right({trees[2138], lumberyards[2138]}), .bottom_left({trees[2186], lumberyards[2186]}), .bottom({trees[2187], lumberyards[2187]}), .bottom_right({trees[2188], lumberyards[2188]}), .init(2'b00), .state({trees[2137], lumberyards[2137]}));
acre acre_42_38 (.clk(clk), .en(en), .top_left({trees[2087], lumberyards[2087]}), .top({trees[2088], lumberyards[2088]}), .top_right({trees[2089], lumberyards[2089]}), .left({trees[2137], lumberyards[2137]}), .right({trees[2139], lumberyards[2139]}), .bottom_left({trees[2187], lumberyards[2187]}), .bottom({trees[2188], lumberyards[2188]}), .bottom_right({trees[2189], lumberyards[2189]}), .init(2'b00), .state({trees[2138], lumberyards[2138]}));
acre acre_42_39 (.clk(clk), .en(en), .top_left({trees[2088], lumberyards[2088]}), .top({trees[2089], lumberyards[2089]}), .top_right({trees[2090], lumberyards[2090]}), .left({trees[2138], lumberyards[2138]}), .right({trees[2140], lumberyards[2140]}), .bottom_left({trees[2188], lumberyards[2188]}), .bottom({trees[2189], lumberyards[2189]}), .bottom_right({trees[2190], lumberyards[2190]}), .init(2'b00), .state({trees[2139], lumberyards[2139]}));
acre acre_42_40 (.clk(clk), .en(en), .top_left({trees[2089], lumberyards[2089]}), .top({trees[2090], lumberyards[2090]}), .top_right({trees[2091], lumberyards[2091]}), .left({trees[2139], lumberyards[2139]}), .right({trees[2141], lumberyards[2141]}), .bottom_left({trees[2189], lumberyards[2189]}), .bottom({trees[2190], lumberyards[2190]}), .bottom_right({trees[2191], lumberyards[2191]}), .init(2'b00), .state({trees[2140], lumberyards[2140]}));
acre acre_42_41 (.clk(clk), .en(en), .top_left({trees[2090], lumberyards[2090]}), .top({trees[2091], lumberyards[2091]}), .top_right({trees[2092], lumberyards[2092]}), .left({trees[2140], lumberyards[2140]}), .right({trees[2142], lumberyards[2142]}), .bottom_left({trees[2190], lumberyards[2190]}), .bottom({trees[2191], lumberyards[2191]}), .bottom_right({trees[2192], lumberyards[2192]}), .init(2'b10), .state({trees[2141], lumberyards[2141]}));
acre acre_42_42 (.clk(clk), .en(en), .top_left({trees[2091], lumberyards[2091]}), .top({trees[2092], lumberyards[2092]}), .top_right({trees[2093], lumberyards[2093]}), .left({trees[2141], lumberyards[2141]}), .right({trees[2143], lumberyards[2143]}), .bottom_left({trees[2191], lumberyards[2191]}), .bottom({trees[2192], lumberyards[2192]}), .bottom_right({trees[2193], lumberyards[2193]}), .init(2'b01), .state({trees[2142], lumberyards[2142]}));
acre acre_42_43 (.clk(clk), .en(en), .top_left({trees[2092], lumberyards[2092]}), .top({trees[2093], lumberyards[2093]}), .top_right({trees[2094], lumberyards[2094]}), .left({trees[2142], lumberyards[2142]}), .right({trees[2144], lumberyards[2144]}), .bottom_left({trees[2192], lumberyards[2192]}), .bottom({trees[2193], lumberyards[2193]}), .bottom_right({trees[2194], lumberyards[2194]}), .init(2'b00), .state({trees[2143], lumberyards[2143]}));
acre acre_42_44 (.clk(clk), .en(en), .top_left({trees[2093], lumberyards[2093]}), .top({trees[2094], lumberyards[2094]}), .top_right({trees[2095], lumberyards[2095]}), .left({trees[2143], lumberyards[2143]}), .right({trees[2145], lumberyards[2145]}), .bottom_left({trees[2193], lumberyards[2193]}), .bottom({trees[2194], lumberyards[2194]}), .bottom_right({trees[2195], lumberyards[2195]}), .init(2'b00), .state({trees[2144], lumberyards[2144]}));
acre acre_42_45 (.clk(clk), .en(en), .top_left({trees[2094], lumberyards[2094]}), .top({trees[2095], lumberyards[2095]}), .top_right({trees[2096], lumberyards[2096]}), .left({trees[2144], lumberyards[2144]}), .right({trees[2146], lumberyards[2146]}), .bottom_left({trees[2194], lumberyards[2194]}), .bottom({trees[2195], lumberyards[2195]}), .bottom_right({trees[2196], lumberyards[2196]}), .init(2'b10), .state({trees[2145], lumberyards[2145]}));
acre acre_42_46 (.clk(clk), .en(en), .top_left({trees[2095], lumberyards[2095]}), .top({trees[2096], lumberyards[2096]}), .top_right({trees[2097], lumberyards[2097]}), .left({trees[2145], lumberyards[2145]}), .right({trees[2147], lumberyards[2147]}), .bottom_left({trees[2195], lumberyards[2195]}), .bottom({trees[2196], lumberyards[2196]}), .bottom_right({trees[2197], lumberyards[2197]}), .init(2'b10), .state({trees[2146], lumberyards[2146]}));
acre acre_42_47 (.clk(clk), .en(en), .top_left({trees[2096], lumberyards[2096]}), .top({trees[2097], lumberyards[2097]}), .top_right({trees[2098], lumberyards[2098]}), .left({trees[2146], lumberyards[2146]}), .right({trees[2148], lumberyards[2148]}), .bottom_left({trees[2196], lumberyards[2196]}), .bottom({trees[2197], lumberyards[2197]}), .bottom_right({trees[2198], lumberyards[2198]}), .init(2'b10), .state({trees[2147], lumberyards[2147]}));
acre acre_42_48 (.clk(clk), .en(en), .top_left({trees[2097], lumberyards[2097]}), .top({trees[2098], lumberyards[2098]}), .top_right({trees[2099], lumberyards[2099]}), .left({trees[2147], lumberyards[2147]}), .right({trees[2149], lumberyards[2149]}), .bottom_left({trees[2197], lumberyards[2197]}), .bottom({trees[2198], lumberyards[2198]}), .bottom_right({trees[2199], lumberyards[2199]}), .init(2'b00), .state({trees[2148], lumberyards[2148]}));
acre acre_42_49 (.clk(clk), .en(en), .top_left({trees[2098], lumberyards[2098]}), .top({trees[2099], lumberyards[2099]}), .top_right(2'b0), .left({trees[2148], lumberyards[2148]}), .right(2'b0), .bottom_left({trees[2198], lumberyards[2198]}), .bottom({trees[2199], lumberyards[2199]}), .bottom_right(2'b0), .init(2'b00), .state({trees[2149], lumberyards[2149]}));
acre acre_43_0 (.clk(clk), .en(en), .top_left(2'b0), .top({trees[2100], lumberyards[2100]}), .top_right({trees[2101], lumberyards[2101]}), .left(2'b0), .right({trees[2151], lumberyards[2151]}), .bottom_left(2'b0), .bottom({trees[2200], lumberyards[2200]}), .bottom_right({trees[2201], lumberyards[2201]}), .init(2'b01), .state({trees[2150], lumberyards[2150]}));
acre acre_43_1 (.clk(clk), .en(en), .top_left({trees[2100], lumberyards[2100]}), .top({trees[2101], lumberyards[2101]}), .top_right({trees[2102], lumberyards[2102]}), .left({trees[2150], lumberyards[2150]}), .right({trees[2152], lumberyards[2152]}), .bottom_left({trees[2200], lumberyards[2200]}), .bottom({trees[2201], lumberyards[2201]}), .bottom_right({trees[2202], lumberyards[2202]}), .init(2'b00), .state({trees[2151], lumberyards[2151]}));
acre acre_43_2 (.clk(clk), .en(en), .top_left({trees[2101], lumberyards[2101]}), .top({trees[2102], lumberyards[2102]}), .top_right({trees[2103], lumberyards[2103]}), .left({trees[2151], lumberyards[2151]}), .right({trees[2153], lumberyards[2153]}), .bottom_left({trees[2201], lumberyards[2201]}), .bottom({trees[2202], lumberyards[2202]}), .bottom_right({trees[2203], lumberyards[2203]}), .init(2'b00), .state({trees[2152], lumberyards[2152]}));
acre acre_43_3 (.clk(clk), .en(en), .top_left({trees[2102], lumberyards[2102]}), .top({trees[2103], lumberyards[2103]}), .top_right({trees[2104], lumberyards[2104]}), .left({trees[2152], lumberyards[2152]}), .right({trees[2154], lumberyards[2154]}), .bottom_left({trees[2202], lumberyards[2202]}), .bottom({trees[2203], lumberyards[2203]}), .bottom_right({trees[2204], lumberyards[2204]}), .init(2'b00), .state({trees[2153], lumberyards[2153]}));
acre acre_43_4 (.clk(clk), .en(en), .top_left({trees[2103], lumberyards[2103]}), .top({trees[2104], lumberyards[2104]}), .top_right({trees[2105], lumberyards[2105]}), .left({trees[2153], lumberyards[2153]}), .right({trees[2155], lumberyards[2155]}), .bottom_left({trees[2203], lumberyards[2203]}), .bottom({trees[2204], lumberyards[2204]}), .bottom_right({trees[2205], lumberyards[2205]}), .init(2'b00), .state({trees[2154], lumberyards[2154]}));
acre acre_43_5 (.clk(clk), .en(en), .top_left({trees[2104], lumberyards[2104]}), .top({trees[2105], lumberyards[2105]}), .top_right({trees[2106], lumberyards[2106]}), .left({trees[2154], lumberyards[2154]}), .right({trees[2156], lumberyards[2156]}), .bottom_left({trees[2204], lumberyards[2204]}), .bottom({trees[2205], lumberyards[2205]}), .bottom_right({trees[2206], lumberyards[2206]}), .init(2'b01), .state({trees[2155], lumberyards[2155]}));
acre acre_43_6 (.clk(clk), .en(en), .top_left({trees[2105], lumberyards[2105]}), .top({trees[2106], lumberyards[2106]}), .top_right({trees[2107], lumberyards[2107]}), .left({trees[2155], lumberyards[2155]}), .right({trees[2157], lumberyards[2157]}), .bottom_left({trees[2205], lumberyards[2205]}), .bottom({trees[2206], lumberyards[2206]}), .bottom_right({trees[2207], lumberyards[2207]}), .init(2'b00), .state({trees[2156], lumberyards[2156]}));
acre acre_43_7 (.clk(clk), .en(en), .top_left({trees[2106], lumberyards[2106]}), .top({trees[2107], lumberyards[2107]}), .top_right({trees[2108], lumberyards[2108]}), .left({trees[2156], lumberyards[2156]}), .right({trees[2158], lumberyards[2158]}), .bottom_left({trees[2206], lumberyards[2206]}), .bottom({trees[2207], lumberyards[2207]}), .bottom_right({trees[2208], lumberyards[2208]}), .init(2'b10), .state({trees[2157], lumberyards[2157]}));
acre acre_43_8 (.clk(clk), .en(en), .top_left({trees[2107], lumberyards[2107]}), .top({trees[2108], lumberyards[2108]}), .top_right({trees[2109], lumberyards[2109]}), .left({trees[2157], lumberyards[2157]}), .right({trees[2159], lumberyards[2159]}), .bottom_left({trees[2207], lumberyards[2207]}), .bottom({trees[2208], lumberyards[2208]}), .bottom_right({trees[2209], lumberyards[2209]}), .init(2'b00), .state({trees[2158], lumberyards[2158]}));
acre acre_43_9 (.clk(clk), .en(en), .top_left({trees[2108], lumberyards[2108]}), .top({trees[2109], lumberyards[2109]}), .top_right({trees[2110], lumberyards[2110]}), .left({trees[2158], lumberyards[2158]}), .right({trees[2160], lumberyards[2160]}), .bottom_left({trees[2208], lumberyards[2208]}), .bottom({trees[2209], lumberyards[2209]}), .bottom_right({trees[2210], lumberyards[2210]}), .init(2'b00), .state({trees[2159], lumberyards[2159]}));
acre acre_43_10 (.clk(clk), .en(en), .top_left({trees[2109], lumberyards[2109]}), .top({trees[2110], lumberyards[2110]}), .top_right({trees[2111], lumberyards[2111]}), .left({trees[2159], lumberyards[2159]}), .right({trees[2161], lumberyards[2161]}), .bottom_left({trees[2209], lumberyards[2209]}), .bottom({trees[2210], lumberyards[2210]}), .bottom_right({trees[2211], lumberyards[2211]}), .init(2'b00), .state({trees[2160], lumberyards[2160]}));
acre acre_43_11 (.clk(clk), .en(en), .top_left({trees[2110], lumberyards[2110]}), .top({trees[2111], lumberyards[2111]}), .top_right({trees[2112], lumberyards[2112]}), .left({trees[2160], lumberyards[2160]}), .right({trees[2162], lumberyards[2162]}), .bottom_left({trees[2210], lumberyards[2210]}), .bottom({trees[2211], lumberyards[2211]}), .bottom_right({trees[2212], lumberyards[2212]}), .init(2'b10), .state({trees[2161], lumberyards[2161]}));
acre acre_43_12 (.clk(clk), .en(en), .top_left({trees[2111], lumberyards[2111]}), .top({trees[2112], lumberyards[2112]}), .top_right({trees[2113], lumberyards[2113]}), .left({trees[2161], lumberyards[2161]}), .right({trees[2163], lumberyards[2163]}), .bottom_left({trees[2211], lumberyards[2211]}), .bottom({trees[2212], lumberyards[2212]}), .bottom_right({trees[2213], lumberyards[2213]}), .init(2'b10), .state({trees[2162], lumberyards[2162]}));
acre acre_43_13 (.clk(clk), .en(en), .top_left({trees[2112], lumberyards[2112]}), .top({trees[2113], lumberyards[2113]}), .top_right({trees[2114], lumberyards[2114]}), .left({trees[2162], lumberyards[2162]}), .right({trees[2164], lumberyards[2164]}), .bottom_left({trees[2212], lumberyards[2212]}), .bottom({trees[2213], lumberyards[2213]}), .bottom_right({trees[2214], lumberyards[2214]}), .init(2'b01), .state({trees[2163], lumberyards[2163]}));
acre acre_43_14 (.clk(clk), .en(en), .top_left({trees[2113], lumberyards[2113]}), .top({trees[2114], lumberyards[2114]}), .top_right({trees[2115], lumberyards[2115]}), .left({trees[2163], lumberyards[2163]}), .right({trees[2165], lumberyards[2165]}), .bottom_left({trees[2213], lumberyards[2213]}), .bottom({trees[2214], lumberyards[2214]}), .bottom_right({trees[2215], lumberyards[2215]}), .init(2'b00), .state({trees[2164], lumberyards[2164]}));
acre acre_43_15 (.clk(clk), .en(en), .top_left({trees[2114], lumberyards[2114]}), .top({trees[2115], lumberyards[2115]}), .top_right({trees[2116], lumberyards[2116]}), .left({trees[2164], lumberyards[2164]}), .right({trees[2166], lumberyards[2166]}), .bottom_left({trees[2214], lumberyards[2214]}), .bottom({trees[2215], lumberyards[2215]}), .bottom_right({trees[2216], lumberyards[2216]}), .init(2'b00), .state({trees[2165], lumberyards[2165]}));
acre acre_43_16 (.clk(clk), .en(en), .top_left({trees[2115], lumberyards[2115]}), .top({trees[2116], lumberyards[2116]}), .top_right({trees[2117], lumberyards[2117]}), .left({trees[2165], lumberyards[2165]}), .right({trees[2167], lumberyards[2167]}), .bottom_left({trees[2215], lumberyards[2215]}), .bottom({trees[2216], lumberyards[2216]}), .bottom_right({trees[2217], lumberyards[2217]}), .init(2'b00), .state({trees[2166], lumberyards[2166]}));
acre acre_43_17 (.clk(clk), .en(en), .top_left({trees[2116], lumberyards[2116]}), .top({trees[2117], lumberyards[2117]}), .top_right({trees[2118], lumberyards[2118]}), .left({trees[2166], lumberyards[2166]}), .right({trees[2168], lumberyards[2168]}), .bottom_left({trees[2216], lumberyards[2216]}), .bottom({trees[2217], lumberyards[2217]}), .bottom_right({trees[2218], lumberyards[2218]}), .init(2'b10), .state({trees[2167], lumberyards[2167]}));
acre acre_43_18 (.clk(clk), .en(en), .top_left({trees[2117], lumberyards[2117]}), .top({trees[2118], lumberyards[2118]}), .top_right({trees[2119], lumberyards[2119]}), .left({trees[2167], lumberyards[2167]}), .right({trees[2169], lumberyards[2169]}), .bottom_left({trees[2217], lumberyards[2217]}), .bottom({trees[2218], lumberyards[2218]}), .bottom_right({trees[2219], lumberyards[2219]}), .init(2'b00), .state({trees[2168], lumberyards[2168]}));
acre acre_43_19 (.clk(clk), .en(en), .top_left({trees[2118], lumberyards[2118]}), .top({trees[2119], lumberyards[2119]}), .top_right({trees[2120], lumberyards[2120]}), .left({trees[2168], lumberyards[2168]}), .right({trees[2170], lumberyards[2170]}), .bottom_left({trees[2218], lumberyards[2218]}), .bottom({trees[2219], lumberyards[2219]}), .bottom_right({trees[2220], lumberyards[2220]}), .init(2'b01), .state({trees[2169], lumberyards[2169]}));
acre acre_43_20 (.clk(clk), .en(en), .top_left({trees[2119], lumberyards[2119]}), .top({trees[2120], lumberyards[2120]}), .top_right({trees[2121], lumberyards[2121]}), .left({trees[2169], lumberyards[2169]}), .right({trees[2171], lumberyards[2171]}), .bottom_left({trees[2219], lumberyards[2219]}), .bottom({trees[2220], lumberyards[2220]}), .bottom_right({trees[2221], lumberyards[2221]}), .init(2'b00), .state({trees[2170], lumberyards[2170]}));
acre acre_43_21 (.clk(clk), .en(en), .top_left({trees[2120], lumberyards[2120]}), .top({trees[2121], lumberyards[2121]}), .top_right({trees[2122], lumberyards[2122]}), .left({trees[2170], lumberyards[2170]}), .right({trees[2172], lumberyards[2172]}), .bottom_left({trees[2220], lumberyards[2220]}), .bottom({trees[2221], lumberyards[2221]}), .bottom_right({trees[2222], lumberyards[2222]}), .init(2'b01), .state({trees[2171], lumberyards[2171]}));
acre acre_43_22 (.clk(clk), .en(en), .top_left({trees[2121], lumberyards[2121]}), .top({trees[2122], lumberyards[2122]}), .top_right({trees[2123], lumberyards[2123]}), .left({trees[2171], lumberyards[2171]}), .right({trees[2173], lumberyards[2173]}), .bottom_left({trees[2221], lumberyards[2221]}), .bottom({trees[2222], lumberyards[2222]}), .bottom_right({trees[2223], lumberyards[2223]}), .init(2'b00), .state({trees[2172], lumberyards[2172]}));
acre acre_43_23 (.clk(clk), .en(en), .top_left({trees[2122], lumberyards[2122]}), .top({trees[2123], lumberyards[2123]}), .top_right({trees[2124], lumberyards[2124]}), .left({trees[2172], lumberyards[2172]}), .right({trees[2174], lumberyards[2174]}), .bottom_left({trees[2222], lumberyards[2222]}), .bottom({trees[2223], lumberyards[2223]}), .bottom_right({trees[2224], lumberyards[2224]}), .init(2'b00), .state({trees[2173], lumberyards[2173]}));
acre acre_43_24 (.clk(clk), .en(en), .top_left({trees[2123], lumberyards[2123]}), .top({trees[2124], lumberyards[2124]}), .top_right({trees[2125], lumberyards[2125]}), .left({trees[2173], lumberyards[2173]}), .right({trees[2175], lumberyards[2175]}), .bottom_left({trees[2223], lumberyards[2223]}), .bottom({trees[2224], lumberyards[2224]}), .bottom_right({trees[2225], lumberyards[2225]}), .init(2'b01), .state({trees[2174], lumberyards[2174]}));
acre acre_43_25 (.clk(clk), .en(en), .top_left({trees[2124], lumberyards[2124]}), .top({trees[2125], lumberyards[2125]}), .top_right({trees[2126], lumberyards[2126]}), .left({trees[2174], lumberyards[2174]}), .right({trees[2176], lumberyards[2176]}), .bottom_left({trees[2224], lumberyards[2224]}), .bottom({trees[2225], lumberyards[2225]}), .bottom_right({trees[2226], lumberyards[2226]}), .init(2'b10), .state({trees[2175], lumberyards[2175]}));
acre acre_43_26 (.clk(clk), .en(en), .top_left({trees[2125], lumberyards[2125]}), .top({trees[2126], lumberyards[2126]}), .top_right({trees[2127], lumberyards[2127]}), .left({trees[2175], lumberyards[2175]}), .right({trees[2177], lumberyards[2177]}), .bottom_left({trees[2225], lumberyards[2225]}), .bottom({trees[2226], lumberyards[2226]}), .bottom_right({trees[2227], lumberyards[2227]}), .init(2'b00), .state({trees[2176], lumberyards[2176]}));
acre acre_43_27 (.clk(clk), .en(en), .top_left({trees[2126], lumberyards[2126]}), .top({trees[2127], lumberyards[2127]}), .top_right({trees[2128], lumberyards[2128]}), .left({trees[2176], lumberyards[2176]}), .right({trees[2178], lumberyards[2178]}), .bottom_left({trees[2226], lumberyards[2226]}), .bottom({trees[2227], lumberyards[2227]}), .bottom_right({trees[2228], lumberyards[2228]}), .init(2'b00), .state({trees[2177], lumberyards[2177]}));
acre acre_43_28 (.clk(clk), .en(en), .top_left({trees[2127], lumberyards[2127]}), .top({trees[2128], lumberyards[2128]}), .top_right({trees[2129], lumberyards[2129]}), .left({trees[2177], lumberyards[2177]}), .right({trees[2179], lumberyards[2179]}), .bottom_left({trees[2227], lumberyards[2227]}), .bottom({trees[2228], lumberyards[2228]}), .bottom_right({trees[2229], lumberyards[2229]}), .init(2'b00), .state({trees[2178], lumberyards[2178]}));
acre acre_43_29 (.clk(clk), .en(en), .top_left({trees[2128], lumberyards[2128]}), .top({trees[2129], lumberyards[2129]}), .top_right({trees[2130], lumberyards[2130]}), .left({trees[2178], lumberyards[2178]}), .right({trees[2180], lumberyards[2180]}), .bottom_left({trees[2228], lumberyards[2228]}), .bottom({trees[2229], lumberyards[2229]}), .bottom_right({trees[2230], lumberyards[2230]}), .init(2'b00), .state({trees[2179], lumberyards[2179]}));
acre acre_43_30 (.clk(clk), .en(en), .top_left({trees[2129], lumberyards[2129]}), .top({trees[2130], lumberyards[2130]}), .top_right({trees[2131], lumberyards[2131]}), .left({trees[2179], lumberyards[2179]}), .right({trees[2181], lumberyards[2181]}), .bottom_left({trees[2229], lumberyards[2229]}), .bottom({trees[2230], lumberyards[2230]}), .bottom_right({trees[2231], lumberyards[2231]}), .init(2'b00), .state({trees[2180], lumberyards[2180]}));
acre acre_43_31 (.clk(clk), .en(en), .top_left({trees[2130], lumberyards[2130]}), .top({trees[2131], lumberyards[2131]}), .top_right({trees[2132], lumberyards[2132]}), .left({trees[2180], lumberyards[2180]}), .right({trees[2182], lumberyards[2182]}), .bottom_left({trees[2230], lumberyards[2230]}), .bottom({trees[2231], lumberyards[2231]}), .bottom_right({trees[2232], lumberyards[2232]}), .init(2'b00), .state({trees[2181], lumberyards[2181]}));
acre acre_43_32 (.clk(clk), .en(en), .top_left({trees[2131], lumberyards[2131]}), .top({trees[2132], lumberyards[2132]}), .top_right({trees[2133], lumberyards[2133]}), .left({trees[2181], lumberyards[2181]}), .right({trees[2183], lumberyards[2183]}), .bottom_left({trees[2231], lumberyards[2231]}), .bottom({trees[2232], lumberyards[2232]}), .bottom_right({trees[2233], lumberyards[2233]}), .init(2'b00), .state({trees[2182], lumberyards[2182]}));
acre acre_43_33 (.clk(clk), .en(en), .top_left({trees[2132], lumberyards[2132]}), .top({trees[2133], lumberyards[2133]}), .top_right({trees[2134], lumberyards[2134]}), .left({trees[2182], lumberyards[2182]}), .right({trees[2184], lumberyards[2184]}), .bottom_left({trees[2232], lumberyards[2232]}), .bottom({trees[2233], lumberyards[2233]}), .bottom_right({trees[2234], lumberyards[2234]}), .init(2'b01), .state({trees[2183], lumberyards[2183]}));
acre acre_43_34 (.clk(clk), .en(en), .top_left({trees[2133], lumberyards[2133]}), .top({trees[2134], lumberyards[2134]}), .top_right({trees[2135], lumberyards[2135]}), .left({trees[2183], lumberyards[2183]}), .right({trees[2185], lumberyards[2185]}), .bottom_left({trees[2233], lumberyards[2233]}), .bottom({trees[2234], lumberyards[2234]}), .bottom_right({trees[2235], lumberyards[2235]}), .init(2'b00), .state({trees[2184], lumberyards[2184]}));
acre acre_43_35 (.clk(clk), .en(en), .top_left({trees[2134], lumberyards[2134]}), .top({trees[2135], lumberyards[2135]}), .top_right({trees[2136], lumberyards[2136]}), .left({trees[2184], lumberyards[2184]}), .right({trees[2186], lumberyards[2186]}), .bottom_left({trees[2234], lumberyards[2234]}), .bottom({trees[2235], lumberyards[2235]}), .bottom_right({trees[2236], lumberyards[2236]}), .init(2'b00), .state({trees[2185], lumberyards[2185]}));
acre acre_43_36 (.clk(clk), .en(en), .top_left({trees[2135], lumberyards[2135]}), .top({trees[2136], lumberyards[2136]}), .top_right({trees[2137], lumberyards[2137]}), .left({trees[2185], lumberyards[2185]}), .right({trees[2187], lumberyards[2187]}), .bottom_left({trees[2235], lumberyards[2235]}), .bottom({trees[2236], lumberyards[2236]}), .bottom_right({trees[2237], lumberyards[2237]}), .init(2'b00), .state({trees[2186], lumberyards[2186]}));
acre acre_43_37 (.clk(clk), .en(en), .top_left({trees[2136], lumberyards[2136]}), .top({trees[2137], lumberyards[2137]}), .top_right({trees[2138], lumberyards[2138]}), .left({trees[2186], lumberyards[2186]}), .right({trees[2188], lumberyards[2188]}), .bottom_left({trees[2236], lumberyards[2236]}), .bottom({trees[2237], lumberyards[2237]}), .bottom_right({trees[2238], lumberyards[2238]}), .init(2'b10), .state({trees[2187], lumberyards[2187]}));
acre acre_43_38 (.clk(clk), .en(en), .top_left({trees[2137], lumberyards[2137]}), .top({trees[2138], lumberyards[2138]}), .top_right({trees[2139], lumberyards[2139]}), .left({trees[2187], lumberyards[2187]}), .right({trees[2189], lumberyards[2189]}), .bottom_left({trees[2237], lumberyards[2237]}), .bottom({trees[2238], lumberyards[2238]}), .bottom_right({trees[2239], lumberyards[2239]}), .init(2'b00), .state({trees[2188], lumberyards[2188]}));
acre acre_43_39 (.clk(clk), .en(en), .top_left({trees[2138], lumberyards[2138]}), .top({trees[2139], lumberyards[2139]}), .top_right({trees[2140], lumberyards[2140]}), .left({trees[2188], lumberyards[2188]}), .right({trees[2190], lumberyards[2190]}), .bottom_left({trees[2238], lumberyards[2238]}), .bottom({trees[2239], lumberyards[2239]}), .bottom_right({trees[2240], lumberyards[2240]}), .init(2'b00), .state({trees[2189], lumberyards[2189]}));
acre acre_43_40 (.clk(clk), .en(en), .top_left({trees[2139], lumberyards[2139]}), .top({trees[2140], lumberyards[2140]}), .top_right({trees[2141], lumberyards[2141]}), .left({trees[2189], lumberyards[2189]}), .right({trees[2191], lumberyards[2191]}), .bottom_left({trees[2239], lumberyards[2239]}), .bottom({trees[2240], lumberyards[2240]}), .bottom_right({trees[2241], lumberyards[2241]}), .init(2'b00), .state({trees[2190], lumberyards[2190]}));
acre acre_43_41 (.clk(clk), .en(en), .top_left({trees[2140], lumberyards[2140]}), .top({trees[2141], lumberyards[2141]}), .top_right({trees[2142], lumberyards[2142]}), .left({trees[2190], lumberyards[2190]}), .right({trees[2192], lumberyards[2192]}), .bottom_left({trees[2240], lumberyards[2240]}), .bottom({trees[2241], lumberyards[2241]}), .bottom_right({trees[2242], lumberyards[2242]}), .init(2'b00), .state({trees[2191], lumberyards[2191]}));
acre acre_43_42 (.clk(clk), .en(en), .top_left({trees[2141], lumberyards[2141]}), .top({trees[2142], lumberyards[2142]}), .top_right({trees[2143], lumberyards[2143]}), .left({trees[2191], lumberyards[2191]}), .right({trees[2193], lumberyards[2193]}), .bottom_left({trees[2241], lumberyards[2241]}), .bottom({trees[2242], lumberyards[2242]}), .bottom_right({trees[2243], lumberyards[2243]}), .init(2'b01), .state({trees[2192], lumberyards[2192]}));
acre acre_43_43 (.clk(clk), .en(en), .top_left({trees[2142], lumberyards[2142]}), .top({trees[2143], lumberyards[2143]}), .top_right({trees[2144], lumberyards[2144]}), .left({trees[2192], lumberyards[2192]}), .right({trees[2194], lumberyards[2194]}), .bottom_left({trees[2242], lumberyards[2242]}), .bottom({trees[2243], lumberyards[2243]}), .bottom_right({trees[2244], lumberyards[2244]}), .init(2'b00), .state({trees[2193], lumberyards[2193]}));
acre acre_43_44 (.clk(clk), .en(en), .top_left({trees[2143], lumberyards[2143]}), .top({trees[2144], lumberyards[2144]}), .top_right({trees[2145], lumberyards[2145]}), .left({trees[2193], lumberyards[2193]}), .right({trees[2195], lumberyards[2195]}), .bottom_left({trees[2243], lumberyards[2243]}), .bottom({trees[2244], lumberyards[2244]}), .bottom_right({trees[2245], lumberyards[2245]}), .init(2'b00), .state({trees[2194], lumberyards[2194]}));
acre acre_43_45 (.clk(clk), .en(en), .top_left({trees[2144], lumberyards[2144]}), .top({trees[2145], lumberyards[2145]}), .top_right({trees[2146], lumberyards[2146]}), .left({trees[2194], lumberyards[2194]}), .right({trees[2196], lumberyards[2196]}), .bottom_left({trees[2244], lumberyards[2244]}), .bottom({trees[2245], lumberyards[2245]}), .bottom_right({trees[2246], lumberyards[2246]}), .init(2'b01), .state({trees[2195], lumberyards[2195]}));
acre acre_43_46 (.clk(clk), .en(en), .top_left({trees[2145], lumberyards[2145]}), .top({trees[2146], lumberyards[2146]}), .top_right({trees[2147], lumberyards[2147]}), .left({trees[2195], lumberyards[2195]}), .right({trees[2197], lumberyards[2197]}), .bottom_left({trees[2245], lumberyards[2245]}), .bottom({trees[2246], lumberyards[2246]}), .bottom_right({trees[2247], lumberyards[2247]}), .init(2'b00), .state({trees[2196], lumberyards[2196]}));
acre acre_43_47 (.clk(clk), .en(en), .top_left({trees[2146], lumberyards[2146]}), .top({trees[2147], lumberyards[2147]}), .top_right({trees[2148], lumberyards[2148]}), .left({trees[2196], lumberyards[2196]}), .right({trees[2198], lumberyards[2198]}), .bottom_left({trees[2246], lumberyards[2246]}), .bottom({trees[2247], lumberyards[2247]}), .bottom_right({trees[2248], lumberyards[2248]}), .init(2'b01), .state({trees[2197], lumberyards[2197]}));
acre acre_43_48 (.clk(clk), .en(en), .top_left({trees[2147], lumberyards[2147]}), .top({trees[2148], lumberyards[2148]}), .top_right({trees[2149], lumberyards[2149]}), .left({trees[2197], lumberyards[2197]}), .right({trees[2199], lumberyards[2199]}), .bottom_left({trees[2247], lumberyards[2247]}), .bottom({trees[2248], lumberyards[2248]}), .bottom_right({trees[2249], lumberyards[2249]}), .init(2'b10), .state({trees[2198], lumberyards[2198]}));
acre acre_43_49 (.clk(clk), .en(en), .top_left({trees[2148], lumberyards[2148]}), .top({trees[2149], lumberyards[2149]}), .top_right(2'b0), .left({trees[2198], lumberyards[2198]}), .right(2'b0), .bottom_left({trees[2248], lumberyards[2248]}), .bottom({trees[2249], lumberyards[2249]}), .bottom_right(2'b0), .init(2'b00), .state({trees[2199], lumberyards[2199]}));
acre acre_44_0 (.clk(clk), .en(en), .top_left(2'b0), .top({trees[2150], lumberyards[2150]}), .top_right({trees[2151], lumberyards[2151]}), .left(2'b0), .right({trees[2201], lumberyards[2201]}), .bottom_left(2'b0), .bottom({trees[2250], lumberyards[2250]}), .bottom_right({trees[2251], lumberyards[2251]}), .init(2'b10), .state({trees[2200], lumberyards[2200]}));
acre acre_44_1 (.clk(clk), .en(en), .top_left({trees[2150], lumberyards[2150]}), .top({trees[2151], lumberyards[2151]}), .top_right({trees[2152], lumberyards[2152]}), .left({trees[2200], lumberyards[2200]}), .right({trees[2202], lumberyards[2202]}), .bottom_left({trees[2250], lumberyards[2250]}), .bottom({trees[2251], lumberyards[2251]}), .bottom_right({trees[2252], lumberyards[2252]}), .init(2'b00), .state({trees[2201], lumberyards[2201]}));
acre acre_44_2 (.clk(clk), .en(en), .top_left({trees[2151], lumberyards[2151]}), .top({trees[2152], lumberyards[2152]}), .top_right({trees[2153], lumberyards[2153]}), .left({trees[2201], lumberyards[2201]}), .right({trees[2203], lumberyards[2203]}), .bottom_left({trees[2251], lumberyards[2251]}), .bottom({trees[2252], lumberyards[2252]}), .bottom_right({trees[2253], lumberyards[2253]}), .init(2'b01), .state({trees[2202], lumberyards[2202]}));
acre acre_44_3 (.clk(clk), .en(en), .top_left({trees[2152], lumberyards[2152]}), .top({trees[2153], lumberyards[2153]}), .top_right({trees[2154], lumberyards[2154]}), .left({trees[2202], lumberyards[2202]}), .right({trees[2204], lumberyards[2204]}), .bottom_left({trees[2252], lumberyards[2252]}), .bottom({trees[2253], lumberyards[2253]}), .bottom_right({trees[2254], lumberyards[2254]}), .init(2'b00), .state({trees[2203], lumberyards[2203]}));
acre acre_44_4 (.clk(clk), .en(en), .top_left({trees[2153], lumberyards[2153]}), .top({trees[2154], lumberyards[2154]}), .top_right({trees[2155], lumberyards[2155]}), .left({trees[2203], lumberyards[2203]}), .right({trees[2205], lumberyards[2205]}), .bottom_left({trees[2253], lumberyards[2253]}), .bottom({trees[2254], lumberyards[2254]}), .bottom_right({trees[2255], lumberyards[2255]}), .init(2'b00), .state({trees[2204], lumberyards[2204]}));
acre acre_44_5 (.clk(clk), .en(en), .top_left({trees[2154], lumberyards[2154]}), .top({trees[2155], lumberyards[2155]}), .top_right({trees[2156], lumberyards[2156]}), .left({trees[2204], lumberyards[2204]}), .right({trees[2206], lumberyards[2206]}), .bottom_left({trees[2254], lumberyards[2254]}), .bottom({trees[2255], lumberyards[2255]}), .bottom_right({trees[2256], lumberyards[2256]}), .init(2'b01), .state({trees[2205], lumberyards[2205]}));
acre acre_44_6 (.clk(clk), .en(en), .top_left({trees[2155], lumberyards[2155]}), .top({trees[2156], lumberyards[2156]}), .top_right({trees[2157], lumberyards[2157]}), .left({trees[2205], lumberyards[2205]}), .right({trees[2207], lumberyards[2207]}), .bottom_left({trees[2255], lumberyards[2255]}), .bottom({trees[2256], lumberyards[2256]}), .bottom_right({trees[2257], lumberyards[2257]}), .init(2'b00), .state({trees[2206], lumberyards[2206]}));
acre acre_44_7 (.clk(clk), .en(en), .top_left({trees[2156], lumberyards[2156]}), .top({trees[2157], lumberyards[2157]}), .top_right({trees[2158], lumberyards[2158]}), .left({trees[2206], lumberyards[2206]}), .right({trees[2208], lumberyards[2208]}), .bottom_left({trees[2256], lumberyards[2256]}), .bottom({trees[2257], lumberyards[2257]}), .bottom_right({trees[2258], lumberyards[2258]}), .init(2'b10), .state({trees[2207], lumberyards[2207]}));
acre acre_44_8 (.clk(clk), .en(en), .top_left({trees[2157], lumberyards[2157]}), .top({trees[2158], lumberyards[2158]}), .top_right({trees[2159], lumberyards[2159]}), .left({trees[2207], lumberyards[2207]}), .right({trees[2209], lumberyards[2209]}), .bottom_left({trees[2257], lumberyards[2257]}), .bottom({trees[2258], lumberyards[2258]}), .bottom_right({trees[2259], lumberyards[2259]}), .init(2'b10), .state({trees[2208], lumberyards[2208]}));
acre acre_44_9 (.clk(clk), .en(en), .top_left({trees[2158], lumberyards[2158]}), .top({trees[2159], lumberyards[2159]}), .top_right({trees[2160], lumberyards[2160]}), .left({trees[2208], lumberyards[2208]}), .right({trees[2210], lumberyards[2210]}), .bottom_left({trees[2258], lumberyards[2258]}), .bottom({trees[2259], lumberyards[2259]}), .bottom_right({trees[2260], lumberyards[2260]}), .init(2'b00), .state({trees[2209], lumberyards[2209]}));
acre acre_44_10 (.clk(clk), .en(en), .top_left({trees[2159], lumberyards[2159]}), .top({trees[2160], lumberyards[2160]}), .top_right({trees[2161], lumberyards[2161]}), .left({trees[2209], lumberyards[2209]}), .right({trees[2211], lumberyards[2211]}), .bottom_left({trees[2259], lumberyards[2259]}), .bottom({trees[2260], lumberyards[2260]}), .bottom_right({trees[2261], lumberyards[2261]}), .init(2'b00), .state({trees[2210], lumberyards[2210]}));
acre acre_44_11 (.clk(clk), .en(en), .top_left({trees[2160], lumberyards[2160]}), .top({trees[2161], lumberyards[2161]}), .top_right({trees[2162], lumberyards[2162]}), .left({trees[2210], lumberyards[2210]}), .right({trees[2212], lumberyards[2212]}), .bottom_left({trees[2260], lumberyards[2260]}), .bottom({trees[2261], lumberyards[2261]}), .bottom_right({trees[2262], lumberyards[2262]}), .init(2'b00), .state({trees[2211], lumberyards[2211]}));
acre acre_44_12 (.clk(clk), .en(en), .top_left({trees[2161], lumberyards[2161]}), .top({trees[2162], lumberyards[2162]}), .top_right({trees[2163], lumberyards[2163]}), .left({trees[2211], lumberyards[2211]}), .right({trees[2213], lumberyards[2213]}), .bottom_left({trees[2261], lumberyards[2261]}), .bottom({trees[2262], lumberyards[2262]}), .bottom_right({trees[2263], lumberyards[2263]}), .init(2'b10), .state({trees[2212], lumberyards[2212]}));
acre acre_44_13 (.clk(clk), .en(en), .top_left({trees[2162], lumberyards[2162]}), .top({trees[2163], lumberyards[2163]}), .top_right({trees[2164], lumberyards[2164]}), .left({trees[2212], lumberyards[2212]}), .right({trees[2214], lumberyards[2214]}), .bottom_left({trees[2262], lumberyards[2262]}), .bottom({trees[2263], lumberyards[2263]}), .bottom_right({trees[2264], lumberyards[2264]}), .init(2'b00), .state({trees[2213], lumberyards[2213]}));
acre acre_44_14 (.clk(clk), .en(en), .top_left({trees[2163], lumberyards[2163]}), .top({trees[2164], lumberyards[2164]}), .top_right({trees[2165], lumberyards[2165]}), .left({trees[2213], lumberyards[2213]}), .right({trees[2215], lumberyards[2215]}), .bottom_left({trees[2263], lumberyards[2263]}), .bottom({trees[2264], lumberyards[2264]}), .bottom_right({trees[2265], lumberyards[2265]}), .init(2'b00), .state({trees[2214], lumberyards[2214]}));
acre acre_44_15 (.clk(clk), .en(en), .top_left({trees[2164], lumberyards[2164]}), .top({trees[2165], lumberyards[2165]}), .top_right({trees[2166], lumberyards[2166]}), .left({trees[2214], lumberyards[2214]}), .right({trees[2216], lumberyards[2216]}), .bottom_left({trees[2264], lumberyards[2264]}), .bottom({trees[2265], lumberyards[2265]}), .bottom_right({trees[2266], lumberyards[2266]}), .init(2'b00), .state({trees[2215], lumberyards[2215]}));
acre acre_44_16 (.clk(clk), .en(en), .top_left({trees[2165], lumberyards[2165]}), .top({trees[2166], lumberyards[2166]}), .top_right({trees[2167], lumberyards[2167]}), .left({trees[2215], lumberyards[2215]}), .right({trees[2217], lumberyards[2217]}), .bottom_left({trees[2265], lumberyards[2265]}), .bottom({trees[2266], lumberyards[2266]}), .bottom_right({trees[2267], lumberyards[2267]}), .init(2'b00), .state({trees[2216], lumberyards[2216]}));
acre acre_44_17 (.clk(clk), .en(en), .top_left({trees[2166], lumberyards[2166]}), .top({trees[2167], lumberyards[2167]}), .top_right({trees[2168], lumberyards[2168]}), .left({trees[2216], lumberyards[2216]}), .right({trees[2218], lumberyards[2218]}), .bottom_left({trees[2266], lumberyards[2266]}), .bottom({trees[2267], lumberyards[2267]}), .bottom_right({trees[2268], lumberyards[2268]}), .init(2'b00), .state({trees[2217], lumberyards[2217]}));
acre acre_44_18 (.clk(clk), .en(en), .top_left({trees[2167], lumberyards[2167]}), .top({trees[2168], lumberyards[2168]}), .top_right({trees[2169], lumberyards[2169]}), .left({trees[2217], lumberyards[2217]}), .right({trees[2219], lumberyards[2219]}), .bottom_left({trees[2267], lumberyards[2267]}), .bottom({trees[2268], lumberyards[2268]}), .bottom_right({trees[2269], lumberyards[2269]}), .init(2'b00), .state({trees[2218], lumberyards[2218]}));
acre acre_44_19 (.clk(clk), .en(en), .top_left({trees[2168], lumberyards[2168]}), .top({trees[2169], lumberyards[2169]}), .top_right({trees[2170], lumberyards[2170]}), .left({trees[2218], lumberyards[2218]}), .right({trees[2220], lumberyards[2220]}), .bottom_left({trees[2268], lumberyards[2268]}), .bottom({trees[2269], lumberyards[2269]}), .bottom_right({trees[2270], lumberyards[2270]}), .init(2'b00), .state({trees[2219], lumberyards[2219]}));
acre acre_44_20 (.clk(clk), .en(en), .top_left({trees[2169], lumberyards[2169]}), .top({trees[2170], lumberyards[2170]}), .top_right({trees[2171], lumberyards[2171]}), .left({trees[2219], lumberyards[2219]}), .right({trees[2221], lumberyards[2221]}), .bottom_left({trees[2269], lumberyards[2269]}), .bottom({trees[2270], lumberyards[2270]}), .bottom_right({trees[2271], lumberyards[2271]}), .init(2'b00), .state({trees[2220], lumberyards[2220]}));
acre acre_44_21 (.clk(clk), .en(en), .top_left({trees[2170], lumberyards[2170]}), .top({trees[2171], lumberyards[2171]}), .top_right({trees[2172], lumberyards[2172]}), .left({trees[2220], lumberyards[2220]}), .right({trees[2222], lumberyards[2222]}), .bottom_left({trees[2270], lumberyards[2270]}), .bottom({trees[2271], lumberyards[2271]}), .bottom_right({trees[2272], lumberyards[2272]}), .init(2'b00), .state({trees[2221], lumberyards[2221]}));
acre acre_44_22 (.clk(clk), .en(en), .top_left({trees[2171], lumberyards[2171]}), .top({trees[2172], lumberyards[2172]}), .top_right({trees[2173], lumberyards[2173]}), .left({trees[2221], lumberyards[2221]}), .right({trees[2223], lumberyards[2223]}), .bottom_left({trees[2271], lumberyards[2271]}), .bottom({trees[2272], lumberyards[2272]}), .bottom_right({trees[2273], lumberyards[2273]}), .init(2'b00), .state({trees[2222], lumberyards[2222]}));
acre acre_44_23 (.clk(clk), .en(en), .top_left({trees[2172], lumberyards[2172]}), .top({trees[2173], lumberyards[2173]}), .top_right({trees[2174], lumberyards[2174]}), .left({trees[2222], lumberyards[2222]}), .right({trees[2224], lumberyards[2224]}), .bottom_left({trees[2272], lumberyards[2272]}), .bottom({trees[2273], lumberyards[2273]}), .bottom_right({trees[2274], lumberyards[2274]}), .init(2'b01), .state({trees[2223], lumberyards[2223]}));
acre acre_44_24 (.clk(clk), .en(en), .top_left({trees[2173], lumberyards[2173]}), .top({trees[2174], lumberyards[2174]}), .top_right({trees[2175], lumberyards[2175]}), .left({trees[2223], lumberyards[2223]}), .right({trees[2225], lumberyards[2225]}), .bottom_left({trees[2273], lumberyards[2273]}), .bottom({trees[2274], lumberyards[2274]}), .bottom_right({trees[2275], lumberyards[2275]}), .init(2'b00), .state({trees[2224], lumberyards[2224]}));
acre acre_44_25 (.clk(clk), .en(en), .top_left({trees[2174], lumberyards[2174]}), .top({trees[2175], lumberyards[2175]}), .top_right({trees[2176], lumberyards[2176]}), .left({trees[2224], lumberyards[2224]}), .right({trees[2226], lumberyards[2226]}), .bottom_left({trees[2274], lumberyards[2274]}), .bottom({trees[2275], lumberyards[2275]}), .bottom_right({trees[2276], lumberyards[2276]}), .init(2'b01), .state({trees[2225], lumberyards[2225]}));
acre acre_44_26 (.clk(clk), .en(en), .top_left({trees[2175], lumberyards[2175]}), .top({trees[2176], lumberyards[2176]}), .top_right({trees[2177], lumberyards[2177]}), .left({trees[2225], lumberyards[2225]}), .right({trees[2227], lumberyards[2227]}), .bottom_left({trees[2275], lumberyards[2275]}), .bottom({trees[2276], lumberyards[2276]}), .bottom_right({trees[2277], lumberyards[2277]}), .init(2'b10), .state({trees[2226], lumberyards[2226]}));
acre acre_44_27 (.clk(clk), .en(en), .top_left({trees[2176], lumberyards[2176]}), .top({trees[2177], lumberyards[2177]}), .top_right({trees[2178], lumberyards[2178]}), .left({trees[2226], lumberyards[2226]}), .right({trees[2228], lumberyards[2228]}), .bottom_left({trees[2276], lumberyards[2276]}), .bottom({trees[2277], lumberyards[2277]}), .bottom_right({trees[2278], lumberyards[2278]}), .init(2'b00), .state({trees[2227], lumberyards[2227]}));
acre acre_44_28 (.clk(clk), .en(en), .top_left({trees[2177], lumberyards[2177]}), .top({trees[2178], lumberyards[2178]}), .top_right({trees[2179], lumberyards[2179]}), .left({trees[2227], lumberyards[2227]}), .right({trees[2229], lumberyards[2229]}), .bottom_left({trees[2277], lumberyards[2277]}), .bottom({trees[2278], lumberyards[2278]}), .bottom_right({trees[2279], lumberyards[2279]}), .init(2'b00), .state({trees[2228], lumberyards[2228]}));
acre acre_44_29 (.clk(clk), .en(en), .top_left({trees[2178], lumberyards[2178]}), .top({trees[2179], lumberyards[2179]}), .top_right({trees[2180], lumberyards[2180]}), .left({trees[2228], lumberyards[2228]}), .right({trees[2230], lumberyards[2230]}), .bottom_left({trees[2278], lumberyards[2278]}), .bottom({trees[2279], lumberyards[2279]}), .bottom_right({trees[2280], lumberyards[2280]}), .init(2'b00), .state({trees[2229], lumberyards[2229]}));
acre acre_44_30 (.clk(clk), .en(en), .top_left({trees[2179], lumberyards[2179]}), .top({trees[2180], lumberyards[2180]}), .top_right({trees[2181], lumberyards[2181]}), .left({trees[2229], lumberyards[2229]}), .right({trees[2231], lumberyards[2231]}), .bottom_left({trees[2279], lumberyards[2279]}), .bottom({trees[2280], lumberyards[2280]}), .bottom_right({trees[2281], lumberyards[2281]}), .init(2'b01), .state({trees[2230], lumberyards[2230]}));
acre acre_44_31 (.clk(clk), .en(en), .top_left({trees[2180], lumberyards[2180]}), .top({trees[2181], lumberyards[2181]}), .top_right({trees[2182], lumberyards[2182]}), .left({trees[2230], lumberyards[2230]}), .right({trees[2232], lumberyards[2232]}), .bottom_left({trees[2280], lumberyards[2280]}), .bottom({trees[2281], lumberyards[2281]}), .bottom_right({trees[2282], lumberyards[2282]}), .init(2'b01), .state({trees[2231], lumberyards[2231]}));
acre acre_44_32 (.clk(clk), .en(en), .top_left({trees[2181], lumberyards[2181]}), .top({trees[2182], lumberyards[2182]}), .top_right({trees[2183], lumberyards[2183]}), .left({trees[2231], lumberyards[2231]}), .right({trees[2233], lumberyards[2233]}), .bottom_left({trees[2281], lumberyards[2281]}), .bottom({trees[2282], lumberyards[2282]}), .bottom_right({trees[2283], lumberyards[2283]}), .init(2'b00), .state({trees[2232], lumberyards[2232]}));
acre acre_44_33 (.clk(clk), .en(en), .top_left({trees[2182], lumberyards[2182]}), .top({trees[2183], lumberyards[2183]}), .top_right({trees[2184], lumberyards[2184]}), .left({trees[2232], lumberyards[2232]}), .right({trees[2234], lumberyards[2234]}), .bottom_left({trees[2282], lumberyards[2282]}), .bottom({trees[2283], lumberyards[2283]}), .bottom_right({trees[2284], lumberyards[2284]}), .init(2'b01), .state({trees[2233], lumberyards[2233]}));
acre acre_44_34 (.clk(clk), .en(en), .top_left({trees[2183], lumberyards[2183]}), .top({trees[2184], lumberyards[2184]}), .top_right({trees[2185], lumberyards[2185]}), .left({trees[2233], lumberyards[2233]}), .right({trees[2235], lumberyards[2235]}), .bottom_left({trees[2283], lumberyards[2283]}), .bottom({trees[2284], lumberyards[2284]}), .bottom_right({trees[2285], lumberyards[2285]}), .init(2'b00), .state({trees[2234], lumberyards[2234]}));
acre acre_44_35 (.clk(clk), .en(en), .top_left({trees[2184], lumberyards[2184]}), .top({trees[2185], lumberyards[2185]}), .top_right({trees[2186], lumberyards[2186]}), .left({trees[2234], lumberyards[2234]}), .right({trees[2236], lumberyards[2236]}), .bottom_left({trees[2284], lumberyards[2284]}), .bottom({trees[2285], lumberyards[2285]}), .bottom_right({trees[2286], lumberyards[2286]}), .init(2'b10), .state({trees[2235], lumberyards[2235]}));
acre acre_44_36 (.clk(clk), .en(en), .top_left({trees[2185], lumberyards[2185]}), .top({trees[2186], lumberyards[2186]}), .top_right({trees[2187], lumberyards[2187]}), .left({trees[2235], lumberyards[2235]}), .right({trees[2237], lumberyards[2237]}), .bottom_left({trees[2285], lumberyards[2285]}), .bottom({trees[2286], lumberyards[2286]}), .bottom_right({trees[2287], lumberyards[2287]}), .init(2'b10), .state({trees[2236], lumberyards[2236]}));
acre acre_44_37 (.clk(clk), .en(en), .top_left({trees[2186], lumberyards[2186]}), .top({trees[2187], lumberyards[2187]}), .top_right({trees[2188], lumberyards[2188]}), .left({trees[2236], lumberyards[2236]}), .right({trees[2238], lumberyards[2238]}), .bottom_left({trees[2286], lumberyards[2286]}), .bottom({trees[2287], lumberyards[2287]}), .bottom_right({trees[2288], lumberyards[2288]}), .init(2'b00), .state({trees[2237], lumberyards[2237]}));
acre acre_44_38 (.clk(clk), .en(en), .top_left({trees[2187], lumberyards[2187]}), .top({trees[2188], lumberyards[2188]}), .top_right({trees[2189], lumberyards[2189]}), .left({trees[2237], lumberyards[2237]}), .right({trees[2239], lumberyards[2239]}), .bottom_left({trees[2287], lumberyards[2287]}), .bottom({trees[2288], lumberyards[2288]}), .bottom_right({trees[2289], lumberyards[2289]}), .init(2'b10), .state({trees[2238], lumberyards[2238]}));
acre acre_44_39 (.clk(clk), .en(en), .top_left({trees[2188], lumberyards[2188]}), .top({trees[2189], lumberyards[2189]}), .top_right({trees[2190], lumberyards[2190]}), .left({trees[2238], lumberyards[2238]}), .right({trees[2240], lumberyards[2240]}), .bottom_left({trees[2288], lumberyards[2288]}), .bottom({trees[2289], lumberyards[2289]}), .bottom_right({trees[2290], lumberyards[2290]}), .init(2'b01), .state({trees[2239], lumberyards[2239]}));
acre acre_44_40 (.clk(clk), .en(en), .top_left({trees[2189], lumberyards[2189]}), .top({trees[2190], lumberyards[2190]}), .top_right({trees[2191], lumberyards[2191]}), .left({trees[2239], lumberyards[2239]}), .right({trees[2241], lumberyards[2241]}), .bottom_left({trees[2289], lumberyards[2289]}), .bottom({trees[2290], lumberyards[2290]}), .bottom_right({trees[2291], lumberyards[2291]}), .init(2'b10), .state({trees[2240], lumberyards[2240]}));
acre acre_44_41 (.clk(clk), .en(en), .top_left({trees[2190], lumberyards[2190]}), .top({trees[2191], lumberyards[2191]}), .top_right({trees[2192], lumberyards[2192]}), .left({trees[2240], lumberyards[2240]}), .right({trees[2242], lumberyards[2242]}), .bottom_left({trees[2290], lumberyards[2290]}), .bottom({trees[2291], lumberyards[2291]}), .bottom_right({trees[2292], lumberyards[2292]}), .init(2'b00), .state({trees[2241], lumberyards[2241]}));
acre acre_44_42 (.clk(clk), .en(en), .top_left({trees[2191], lumberyards[2191]}), .top({trees[2192], lumberyards[2192]}), .top_right({trees[2193], lumberyards[2193]}), .left({trees[2241], lumberyards[2241]}), .right({trees[2243], lumberyards[2243]}), .bottom_left({trees[2291], lumberyards[2291]}), .bottom({trees[2292], lumberyards[2292]}), .bottom_right({trees[2293], lumberyards[2293]}), .init(2'b00), .state({trees[2242], lumberyards[2242]}));
acre acre_44_43 (.clk(clk), .en(en), .top_left({trees[2192], lumberyards[2192]}), .top({trees[2193], lumberyards[2193]}), .top_right({trees[2194], lumberyards[2194]}), .left({trees[2242], lumberyards[2242]}), .right({trees[2244], lumberyards[2244]}), .bottom_left({trees[2292], lumberyards[2292]}), .bottom({trees[2293], lumberyards[2293]}), .bottom_right({trees[2294], lumberyards[2294]}), .init(2'b00), .state({trees[2243], lumberyards[2243]}));
acre acre_44_44 (.clk(clk), .en(en), .top_left({trees[2193], lumberyards[2193]}), .top({trees[2194], lumberyards[2194]}), .top_right({trees[2195], lumberyards[2195]}), .left({trees[2243], lumberyards[2243]}), .right({trees[2245], lumberyards[2245]}), .bottom_left({trees[2293], lumberyards[2293]}), .bottom({trees[2294], lumberyards[2294]}), .bottom_right({trees[2295], lumberyards[2295]}), .init(2'b00), .state({trees[2244], lumberyards[2244]}));
acre acre_44_45 (.clk(clk), .en(en), .top_left({trees[2194], lumberyards[2194]}), .top({trees[2195], lumberyards[2195]}), .top_right({trees[2196], lumberyards[2196]}), .left({trees[2244], lumberyards[2244]}), .right({trees[2246], lumberyards[2246]}), .bottom_left({trees[2294], lumberyards[2294]}), .bottom({trees[2295], lumberyards[2295]}), .bottom_right({trees[2296], lumberyards[2296]}), .init(2'b00), .state({trees[2245], lumberyards[2245]}));
acre acre_44_46 (.clk(clk), .en(en), .top_left({trees[2195], lumberyards[2195]}), .top({trees[2196], lumberyards[2196]}), .top_right({trees[2197], lumberyards[2197]}), .left({trees[2245], lumberyards[2245]}), .right({trees[2247], lumberyards[2247]}), .bottom_left({trees[2295], lumberyards[2295]}), .bottom({trees[2296], lumberyards[2296]}), .bottom_right({trees[2297], lumberyards[2297]}), .init(2'b00), .state({trees[2246], lumberyards[2246]}));
acre acre_44_47 (.clk(clk), .en(en), .top_left({trees[2196], lumberyards[2196]}), .top({trees[2197], lumberyards[2197]}), .top_right({trees[2198], lumberyards[2198]}), .left({trees[2246], lumberyards[2246]}), .right({trees[2248], lumberyards[2248]}), .bottom_left({trees[2296], lumberyards[2296]}), .bottom({trees[2297], lumberyards[2297]}), .bottom_right({trees[2298], lumberyards[2298]}), .init(2'b00), .state({trees[2247], lumberyards[2247]}));
acre acre_44_48 (.clk(clk), .en(en), .top_left({trees[2197], lumberyards[2197]}), .top({trees[2198], lumberyards[2198]}), .top_right({trees[2199], lumberyards[2199]}), .left({trees[2247], lumberyards[2247]}), .right({trees[2249], lumberyards[2249]}), .bottom_left({trees[2297], lumberyards[2297]}), .bottom({trees[2298], lumberyards[2298]}), .bottom_right({trees[2299], lumberyards[2299]}), .init(2'b00), .state({trees[2248], lumberyards[2248]}));
acre acre_44_49 (.clk(clk), .en(en), .top_left({trees[2198], lumberyards[2198]}), .top({trees[2199], lumberyards[2199]}), .top_right(2'b0), .left({trees[2248], lumberyards[2248]}), .right(2'b0), .bottom_left({trees[2298], lumberyards[2298]}), .bottom({trees[2299], lumberyards[2299]}), .bottom_right(2'b0), .init(2'b00), .state({trees[2249], lumberyards[2249]}));
acre acre_45_0 (.clk(clk), .en(en), .top_left(2'b0), .top({trees[2200], lumberyards[2200]}), .top_right({trees[2201], lumberyards[2201]}), .left(2'b0), .right({trees[2251], lumberyards[2251]}), .bottom_left(2'b0), .bottom({trees[2300], lumberyards[2300]}), .bottom_right({trees[2301], lumberyards[2301]}), .init(2'b00), .state({trees[2250], lumberyards[2250]}));
acre acre_45_1 (.clk(clk), .en(en), .top_left({trees[2200], lumberyards[2200]}), .top({trees[2201], lumberyards[2201]}), .top_right({trees[2202], lumberyards[2202]}), .left({trees[2250], lumberyards[2250]}), .right({trees[2252], lumberyards[2252]}), .bottom_left({trees[2300], lumberyards[2300]}), .bottom({trees[2301], lumberyards[2301]}), .bottom_right({trees[2302], lumberyards[2302]}), .init(2'b00), .state({trees[2251], lumberyards[2251]}));
acre acre_45_2 (.clk(clk), .en(en), .top_left({trees[2201], lumberyards[2201]}), .top({trees[2202], lumberyards[2202]}), .top_right({trees[2203], lumberyards[2203]}), .left({trees[2251], lumberyards[2251]}), .right({trees[2253], lumberyards[2253]}), .bottom_left({trees[2301], lumberyards[2301]}), .bottom({trees[2302], lumberyards[2302]}), .bottom_right({trees[2303], lumberyards[2303]}), .init(2'b01), .state({trees[2252], lumberyards[2252]}));
acre acre_45_3 (.clk(clk), .en(en), .top_left({trees[2202], lumberyards[2202]}), .top({trees[2203], lumberyards[2203]}), .top_right({trees[2204], lumberyards[2204]}), .left({trees[2252], lumberyards[2252]}), .right({trees[2254], lumberyards[2254]}), .bottom_left({trees[2302], lumberyards[2302]}), .bottom({trees[2303], lumberyards[2303]}), .bottom_right({trees[2304], lumberyards[2304]}), .init(2'b00), .state({trees[2253], lumberyards[2253]}));
acre acre_45_4 (.clk(clk), .en(en), .top_left({trees[2203], lumberyards[2203]}), .top({trees[2204], lumberyards[2204]}), .top_right({trees[2205], lumberyards[2205]}), .left({trees[2253], lumberyards[2253]}), .right({trees[2255], lumberyards[2255]}), .bottom_left({trees[2303], lumberyards[2303]}), .bottom({trees[2304], lumberyards[2304]}), .bottom_right({trees[2305], lumberyards[2305]}), .init(2'b01), .state({trees[2254], lumberyards[2254]}));
acre acre_45_5 (.clk(clk), .en(en), .top_left({trees[2204], lumberyards[2204]}), .top({trees[2205], lumberyards[2205]}), .top_right({trees[2206], lumberyards[2206]}), .left({trees[2254], lumberyards[2254]}), .right({trees[2256], lumberyards[2256]}), .bottom_left({trees[2304], lumberyards[2304]}), .bottom({trees[2305], lumberyards[2305]}), .bottom_right({trees[2306], lumberyards[2306]}), .init(2'b01), .state({trees[2255], lumberyards[2255]}));
acre acre_45_6 (.clk(clk), .en(en), .top_left({trees[2205], lumberyards[2205]}), .top({trees[2206], lumberyards[2206]}), .top_right({trees[2207], lumberyards[2207]}), .left({trees[2255], lumberyards[2255]}), .right({trees[2257], lumberyards[2257]}), .bottom_left({trees[2305], lumberyards[2305]}), .bottom({trees[2306], lumberyards[2306]}), .bottom_right({trees[2307], lumberyards[2307]}), .init(2'b10), .state({trees[2256], lumberyards[2256]}));
acre acre_45_7 (.clk(clk), .en(en), .top_left({trees[2206], lumberyards[2206]}), .top({trees[2207], lumberyards[2207]}), .top_right({trees[2208], lumberyards[2208]}), .left({trees[2256], lumberyards[2256]}), .right({trees[2258], lumberyards[2258]}), .bottom_left({trees[2306], lumberyards[2306]}), .bottom({trees[2307], lumberyards[2307]}), .bottom_right({trees[2308], lumberyards[2308]}), .init(2'b01), .state({trees[2257], lumberyards[2257]}));
acre acre_45_8 (.clk(clk), .en(en), .top_left({trees[2207], lumberyards[2207]}), .top({trees[2208], lumberyards[2208]}), .top_right({trees[2209], lumberyards[2209]}), .left({trees[2257], lumberyards[2257]}), .right({trees[2259], lumberyards[2259]}), .bottom_left({trees[2307], lumberyards[2307]}), .bottom({trees[2308], lumberyards[2308]}), .bottom_right({trees[2309], lumberyards[2309]}), .init(2'b01), .state({trees[2258], lumberyards[2258]}));
acre acre_45_9 (.clk(clk), .en(en), .top_left({trees[2208], lumberyards[2208]}), .top({trees[2209], lumberyards[2209]}), .top_right({trees[2210], lumberyards[2210]}), .left({trees[2258], lumberyards[2258]}), .right({trees[2260], lumberyards[2260]}), .bottom_left({trees[2308], lumberyards[2308]}), .bottom({trees[2309], lumberyards[2309]}), .bottom_right({trees[2310], lumberyards[2310]}), .init(2'b00), .state({trees[2259], lumberyards[2259]}));
acre acre_45_10 (.clk(clk), .en(en), .top_left({trees[2209], lumberyards[2209]}), .top({trees[2210], lumberyards[2210]}), .top_right({trees[2211], lumberyards[2211]}), .left({trees[2259], lumberyards[2259]}), .right({trees[2261], lumberyards[2261]}), .bottom_left({trees[2309], lumberyards[2309]}), .bottom({trees[2310], lumberyards[2310]}), .bottom_right({trees[2311], lumberyards[2311]}), .init(2'b00), .state({trees[2260], lumberyards[2260]}));
acre acre_45_11 (.clk(clk), .en(en), .top_left({trees[2210], lumberyards[2210]}), .top({trees[2211], lumberyards[2211]}), .top_right({trees[2212], lumberyards[2212]}), .left({trees[2260], lumberyards[2260]}), .right({trees[2262], lumberyards[2262]}), .bottom_left({trees[2310], lumberyards[2310]}), .bottom({trees[2311], lumberyards[2311]}), .bottom_right({trees[2312], lumberyards[2312]}), .init(2'b10), .state({trees[2261], lumberyards[2261]}));
acre acre_45_12 (.clk(clk), .en(en), .top_left({trees[2211], lumberyards[2211]}), .top({trees[2212], lumberyards[2212]}), .top_right({trees[2213], lumberyards[2213]}), .left({trees[2261], lumberyards[2261]}), .right({trees[2263], lumberyards[2263]}), .bottom_left({trees[2311], lumberyards[2311]}), .bottom({trees[2312], lumberyards[2312]}), .bottom_right({trees[2313], lumberyards[2313]}), .init(2'b00), .state({trees[2262], lumberyards[2262]}));
acre acre_45_13 (.clk(clk), .en(en), .top_left({trees[2212], lumberyards[2212]}), .top({trees[2213], lumberyards[2213]}), .top_right({trees[2214], lumberyards[2214]}), .left({trees[2262], lumberyards[2262]}), .right({trees[2264], lumberyards[2264]}), .bottom_left({trees[2312], lumberyards[2312]}), .bottom({trees[2313], lumberyards[2313]}), .bottom_right({trees[2314], lumberyards[2314]}), .init(2'b01), .state({trees[2263], lumberyards[2263]}));
acre acre_45_14 (.clk(clk), .en(en), .top_left({trees[2213], lumberyards[2213]}), .top({trees[2214], lumberyards[2214]}), .top_right({trees[2215], lumberyards[2215]}), .left({trees[2263], lumberyards[2263]}), .right({trees[2265], lumberyards[2265]}), .bottom_left({trees[2313], lumberyards[2313]}), .bottom({trees[2314], lumberyards[2314]}), .bottom_right({trees[2315], lumberyards[2315]}), .init(2'b10), .state({trees[2264], lumberyards[2264]}));
acre acre_45_15 (.clk(clk), .en(en), .top_left({trees[2214], lumberyards[2214]}), .top({trees[2215], lumberyards[2215]}), .top_right({trees[2216], lumberyards[2216]}), .left({trees[2264], lumberyards[2264]}), .right({trees[2266], lumberyards[2266]}), .bottom_left({trees[2314], lumberyards[2314]}), .bottom({trees[2315], lumberyards[2315]}), .bottom_right({trees[2316], lumberyards[2316]}), .init(2'b00), .state({trees[2265], lumberyards[2265]}));
acre acre_45_16 (.clk(clk), .en(en), .top_left({trees[2215], lumberyards[2215]}), .top({trees[2216], lumberyards[2216]}), .top_right({trees[2217], lumberyards[2217]}), .left({trees[2265], lumberyards[2265]}), .right({trees[2267], lumberyards[2267]}), .bottom_left({trees[2315], lumberyards[2315]}), .bottom({trees[2316], lumberyards[2316]}), .bottom_right({trees[2317], lumberyards[2317]}), .init(2'b01), .state({trees[2266], lumberyards[2266]}));
acre acre_45_17 (.clk(clk), .en(en), .top_left({trees[2216], lumberyards[2216]}), .top({trees[2217], lumberyards[2217]}), .top_right({trees[2218], lumberyards[2218]}), .left({trees[2266], lumberyards[2266]}), .right({trees[2268], lumberyards[2268]}), .bottom_left({trees[2316], lumberyards[2316]}), .bottom({trees[2317], lumberyards[2317]}), .bottom_right({trees[2318], lumberyards[2318]}), .init(2'b01), .state({trees[2267], lumberyards[2267]}));
acre acre_45_18 (.clk(clk), .en(en), .top_left({trees[2217], lumberyards[2217]}), .top({trees[2218], lumberyards[2218]}), .top_right({trees[2219], lumberyards[2219]}), .left({trees[2267], lumberyards[2267]}), .right({trees[2269], lumberyards[2269]}), .bottom_left({trees[2317], lumberyards[2317]}), .bottom({trees[2318], lumberyards[2318]}), .bottom_right({trees[2319], lumberyards[2319]}), .init(2'b00), .state({trees[2268], lumberyards[2268]}));
acre acre_45_19 (.clk(clk), .en(en), .top_left({trees[2218], lumberyards[2218]}), .top({trees[2219], lumberyards[2219]}), .top_right({trees[2220], lumberyards[2220]}), .left({trees[2268], lumberyards[2268]}), .right({trees[2270], lumberyards[2270]}), .bottom_left({trees[2318], lumberyards[2318]}), .bottom({trees[2319], lumberyards[2319]}), .bottom_right({trees[2320], lumberyards[2320]}), .init(2'b10), .state({trees[2269], lumberyards[2269]}));
acre acre_45_20 (.clk(clk), .en(en), .top_left({trees[2219], lumberyards[2219]}), .top({trees[2220], lumberyards[2220]}), .top_right({trees[2221], lumberyards[2221]}), .left({trees[2269], lumberyards[2269]}), .right({trees[2271], lumberyards[2271]}), .bottom_left({trees[2319], lumberyards[2319]}), .bottom({trees[2320], lumberyards[2320]}), .bottom_right({trees[2321], lumberyards[2321]}), .init(2'b00), .state({trees[2270], lumberyards[2270]}));
acre acre_45_21 (.clk(clk), .en(en), .top_left({trees[2220], lumberyards[2220]}), .top({trees[2221], lumberyards[2221]}), .top_right({trees[2222], lumberyards[2222]}), .left({trees[2270], lumberyards[2270]}), .right({trees[2272], lumberyards[2272]}), .bottom_left({trees[2320], lumberyards[2320]}), .bottom({trees[2321], lumberyards[2321]}), .bottom_right({trees[2322], lumberyards[2322]}), .init(2'b00), .state({trees[2271], lumberyards[2271]}));
acre acre_45_22 (.clk(clk), .en(en), .top_left({trees[2221], lumberyards[2221]}), .top({trees[2222], lumberyards[2222]}), .top_right({trees[2223], lumberyards[2223]}), .left({trees[2271], lumberyards[2271]}), .right({trees[2273], lumberyards[2273]}), .bottom_left({trees[2321], lumberyards[2321]}), .bottom({trees[2322], lumberyards[2322]}), .bottom_right({trees[2323], lumberyards[2323]}), .init(2'b00), .state({trees[2272], lumberyards[2272]}));
acre acre_45_23 (.clk(clk), .en(en), .top_left({trees[2222], lumberyards[2222]}), .top({trees[2223], lumberyards[2223]}), .top_right({trees[2224], lumberyards[2224]}), .left({trees[2272], lumberyards[2272]}), .right({trees[2274], lumberyards[2274]}), .bottom_left({trees[2322], lumberyards[2322]}), .bottom({trees[2323], lumberyards[2323]}), .bottom_right({trees[2324], lumberyards[2324]}), .init(2'b00), .state({trees[2273], lumberyards[2273]}));
acre acre_45_24 (.clk(clk), .en(en), .top_left({trees[2223], lumberyards[2223]}), .top({trees[2224], lumberyards[2224]}), .top_right({trees[2225], lumberyards[2225]}), .left({trees[2273], lumberyards[2273]}), .right({trees[2275], lumberyards[2275]}), .bottom_left({trees[2323], lumberyards[2323]}), .bottom({trees[2324], lumberyards[2324]}), .bottom_right({trees[2325], lumberyards[2325]}), .init(2'b00), .state({trees[2274], lumberyards[2274]}));
acre acre_45_25 (.clk(clk), .en(en), .top_left({trees[2224], lumberyards[2224]}), .top({trees[2225], lumberyards[2225]}), .top_right({trees[2226], lumberyards[2226]}), .left({trees[2274], lumberyards[2274]}), .right({trees[2276], lumberyards[2276]}), .bottom_left({trees[2324], lumberyards[2324]}), .bottom({trees[2325], lumberyards[2325]}), .bottom_right({trees[2326], lumberyards[2326]}), .init(2'b01), .state({trees[2275], lumberyards[2275]}));
acre acre_45_26 (.clk(clk), .en(en), .top_left({trees[2225], lumberyards[2225]}), .top({trees[2226], lumberyards[2226]}), .top_right({trees[2227], lumberyards[2227]}), .left({trees[2275], lumberyards[2275]}), .right({trees[2277], lumberyards[2277]}), .bottom_left({trees[2325], lumberyards[2325]}), .bottom({trees[2326], lumberyards[2326]}), .bottom_right({trees[2327], lumberyards[2327]}), .init(2'b00), .state({trees[2276], lumberyards[2276]}));
acre acre_45_27 (.clk(clk), .en(en), .top_left({trees[2226], lumberyards[2226]}), .top({trees[2227], lumberyards[2227]}), .top_right({trees[2228], lumberyards[2228]}), .left({trees[2276], lumberyards[2276]}), .right({trees[2278], lumberyards[2278]}), .bottom_left({trees[2326], lumberyards[2326]}), .bottom({trees[2327], lumberyards[2327]}), .bottom_right({trees[2328], lumberyards[2328]}), .init(2'b00), .state({trees[2277], lumberyards[2277]}));
acre acre_45_28 (.clk(clk), .en(en), .top_left({trees[2227], lumberyards[2227]}), .top({trees[2228], lumberyards[2228]}), .top_right({trees[2229], lumberyards[2229]}), .left({trees[2277], lumberyards[2277]}), .right({trees[2279], lumberyards[2279]}), .bottom_left({trees[2327], lumberyards[2327]}), .bottom({trees[2328], lumberyards[2328]}), .bottom_right({trees[2329], lumberyards[2329]}), .init(2'b00), .state({trees[2278], lumberyards[2278]}));
acre acre_45_29 (.clk(clk), .en(en), .top_left({trees[2228], lumberyards[2228]}), .top({trees[2229], lumberyards[2229]}), .top_right({trees[2230], lumberyards[2230]}), .left({trees[2278], lumberyards[2278]}), .right({trees[2280], lumberyards[2280]}), .bottom_left({trees[2328], lumberyards[2328]}), .bottom({trees[2329], lumberyards[2329]}), .bottom_right({trees[2330], lumberyards[2330]}), .init(2'b00), .state({trees[2279], lumberyards[2279]}));
acre acre_45_30 (.clk(clk), .en(en), .top_left({trees[2229], lumberyards[2229]}), .top({trees[2230], lumberyards[2230]}), .top_right({trees[2231], lumberyards[2231]}), .left({trees[2279], lumberyards[2279]}), .right({trees[2281], lumberyards[2281]}), .bottom_left({trees[2329], lumberyards[2329]}), .bottom({trees[2330], lumberyards[2330]}), .bottom_right({trees[2331], lumberyards[2331]}), .init(2'b01), .state({trees[2280], lumberyards[2280]}));
acre acre_45_31 (.clk(clk), .en(en), .top_left({trees[2230], lumberyards[2230]}), .top({trees[2231], lumberyards[2231]}), .top_right({trees[2232], lumberyards[2232]}), .left({trees[2280], lumberyards[2280]}), .right({trees[2282], lumberyards[2282]}), .bottom_left({trees[2330], lumberyards[2330]}), .bottom({trees[2331], lumberyards[2331]}), .bottom_right({trees[2332], lumberyards[2332]}), .init(2'b00), .state({trees[2281], lumberyards[2281]}));
acre acre_45_32 (.clk(clk), .en(en), .top_left({trees[2231], lumberyards[2231]}), .top({trees[2232], lumberyards[2232]}), .top_right({trees[2233], lumberyards[2233]}), .left({trees[2281], lumberyards[2281]}), .right({trees[2283], lumberyards[2283]}), .bottom_left({trees[2331], lumberyards[2331]}), .bottom({trees[2332], lumberyards[2332]}), .bottom_right({trees[2333], lumberyards[2333]}), .init(2'b00), .state({trees[2282], lumberyards[2282]}));
acre acre_45_33 (.clk(clk), .en(en), .top_left({trees[2232], lumberyards[2232]}), .top({trees[2233], lumberyards[2233]}), .top_right({trees[2234], lumberyards[2234]}), .left({trees[2282], lumberyards[2282]}), .right({trees[2284], lumberyards[2284]}), .bottom_left({trees[2332], lumberyards[2332]}), .bottom({trees[2333], lumberyards[2333]}), .bottom_right({trees[2334], lumberyards[2334]}), .init(2'b00), .state({trees[2283], lumberyards[2283]}));
acre acre_45_34 (.clk(clk), .en(en), .top_left({trees[2233], lumberyards[2233]}), .top({trees[2234], lumberyards[2234]}), .top_right({trees[2235], lumberyards[2235]}), .left({trees[2283], lumberyards[2283]}), .right({trees[2285], lumberyards[2285]}), .bottom_left({trees[2333], lumberyards[2333]}), .bottom({trees[2334], lumberyards[2334]}), .bottom_right({trees[2335], lumberyards[2335]}), .init(2'b10), .state({trees[2284], lumberyards[2284]}));
acre acre_45_35 (.clk(clk), .en(en), .top_left({trees[2234], lumberyards[2234]}), .top({trees[2235], lumberyards[2235]}), .top_right({trees[2236], lumberyards[2236]}), .left({trees[2284], lumberyards[2284]}), .right({trees[2286], lumberyards[2286]}), .bottom_left({trees[2334], lumberyards[2334]}), .bottom({trees[2335], lumberyards[2335]}), .bottom_right({trees[2336], lumberyards[2336]}), .init(2'b00), .state({trees[2285], lumberyards[2285]}));
acre acre_45_36 (.clk(clk), .en(en), .top_left({trees[2235], lumberyards[2235]}), .top({trees[2236], lumberyards[2236]}), .top_right({trees[2237], lumberyards[2237]}), .left({trees[2285], lumberyards[2285]}), .right({trees[2287], lumberyards[2287]}), .bottom_left({trees[2335], lumberyards[2335]}), .bottom({trees[2336], lumberyards[2336]}), .bottom_right({trees[2337], lumberyards[2337]}), .init(2'b10), .state({trees[2286], lumberyards[2286]}));
acre acre_45_37 (.clk(clk), .en(en), .top_left({trees[2236], lumberyards[2236]}), .top({trees[2237], lumberyards[2237]}), .top_right({trees[2238], lumberyards[2238]}), .left({trees[2286], lumberyards[2286]}), .right({trees[2288], lumberyards[2288]}), .bottom_left({trees[2336], lumberyards[2336]}), .bottom({trees[2337], lumberyards[2337]}), .bottom_right({trees[2338], lumberyards[2338]}), .init(2'b01), .state({trees[2287], lumberyards[2287]}));
acre acre_45_38 (.clk(clk), .en(en), .top_left({trees[2237], lumberyards[2237]}), .top({trees[2238], lumberyards[2238]}), .top_right({trees[2239], lumberyards[2239]}), .left({trees[2287], lumberyards[2287]}), .right({trees[2289], lumberyards[2289]}), .bottom_left({trees[2337], lumberyards[2337]}), .bottom({trees[2338], lumberyards[2338]}), .bottom_right({trees[2339], lumberyards[2339]}), .init(2'b01), .state({trees[2288], lumberyards[2288]}));
acre acre_45_39 (.clk(clk), .en(en), .top_left({trees[2238], lumberyards[2238]}), .top({trees[2239], lumberyards[2239]}), .top_right({trees[2240], lumberyards[2240]}), .left({trees[2288], lumberyards[2288]}), .right({trees[2290], lumberyards[2290]}), .bottom_left({trees[2338], lumberyards[2338]}), .bottom({trees[2339], lumberyards[2339]}), .bottom_right({trees[2340], lumberyards[2340]}), .init(2'b00), .state({trees[2289], lumberyards[2289]}));
acre acre_45_40 (.clk(clk), .en(en), .top_left({trees[2239], lumberyards[2239]}), .top({trees[2240], lumberyards[2240]}), .top_right({trees[2241], lumberyards[2241]}), .left({trees[2289], lumberyards[2289]}), .right({trees[2291], lumberyards[2291]}), .bottom_left({trees[2339], lumberyards[2339]}), .bottom({trees[2340], lumberyards[2340]}), .bottom_right({trees[2341], lumberyards[2341]}), .init(2'b00), .state({trees[2290], lumberyards[2290]}));
acre acre_45_41 (.clk(clk), .en(en), .top_left({trees[2240], lumberyards[2240]}), .top({trees[2241], lumberyards[2241]}), .top_right({trees[2242], lumberyards[2242]}), .left({trees[2290], lumberyards[2290]}), .right({trees[2292], lumberyards[2292]}), .bottom_left({trees[2340], lumberyards[2340]}), .bottom({trees[2341], lumberyards[2341]}), .bottom_right({trees[2342], lumberyards[2342]}), .init(2'b00), .state({trees[2291], lumberyards[2291]}));
acre acre_45_42 (.clk(clk), .en(en), .top_left({trees[2241], lumberyards[2241]}), .top({trees[2242], lumberyards[2242]}), .top_right({trees[2243], lumberyards[2243]}), .left({trees[2291], lumberyards[2291]}), .right({trees[2293], lumberyards[2293]}), .bottom_left({trees[2341], lumberyards[2341]}), .bottom({trees[2342], lumberyards[2342]}), .bottom_right({trees[2343], lumberyards[2343]}), .init(2'b00), .state({trees[2292], lumberyards[2292]}));
acre acre_45_43 (.clk(clk), .en(en), .top_left({trees[2242], lumberyards[2242]}), .top({trees[2243], lumberyards[2243]}), .top_right({trees[2244], lumberyards[2244]}), .left({trees[2292], lumberyards[2292]}), .right({trees[2294], lumberyards[2294]}), .bottom_left({trees[2342], lumberyards[2342]}), .bottom({trees[2343], lumberyards[2343]}), .bottom_right({trees[2344], lumberyards[2344]}), .init(2'b10), .state({trees[2293], lumberyards[2293]}));
acre acre_45_44 (.clk(clk), .en(en), .top_left({trees[2243], lumberyards[2243]}), .top({trees[2244], lumberyards[2244]}), .top_right({trees[2245], lumberyards[2245]}), .left({trees[2293], lumberyards[2293]}), .right({trees[2295], lumberyards[2295]}), .bottom_left({trees[2343], lumberyards[2343]}), .bottom({trees[2344], lumberyards[2344]}), .bottom_right({trees[2345], lumberyards[2345]}), .init(2'b00), .state({trees[2294], lumberyards[2294]}));
acre acre_45_45 (.clk(clk), .en(en), .top_left({trees[2244], lumberyards[2244]}), .top({trees[2245], lumberyards[2245]}), .top_right({trees[2246], lumberyards[2246]}), .left({trees[2294], lumberyards[2294]}), .right({trees[2296], lumberyards[2296]}), .bottom_left({trees[2344], lumberyards[2344]}), .bottom({trees[2345], lumberyards[2345]}), .bottom_right({trees[2346], lumberyards[2346]}), .init(2'b00), .state({trees[2295], lumberyards[2295]}));
acre acre_45_46 (.clk(clk), .en(en), .top_left({trees[2245], lumberyards[2245]}), .top({trees[2246], lumberyards[2246]}), .top_right({trees[2247], lumberyards[2247]}), .left({trees[2295], lumberyards[2295]}), .right({trees[2297], lumberyards[2297]}), .bottom_left({trees[2345], lumberyards[2345]}), .bottom({trees[2346], lumberyards[2346]}), .bottom_right({trees[2347], lumberyards[2347]}), .init(2'b00), .state({trees[2296], lumberyards[2296]}));
acre acre_45_47 (.clk(clk), .en(en), .top_left({trees[2246], lumberyards[2246]}), .top({trees[2247], lumberyards[2247]}), .top_right({trees[2248], lumberyards[2248]}), .left({trees[2296], lumberyards[2296]}), .right({trees[2298], lumberyards[2298]}), .bottom_left({trees[2346], lumberyards[2346]}), .bottom({trees[2347], lumberyards[2347]}), .bottom_right({trees[2348], lumberyards[2348]}), .init(2'b00), .state({trees[2297], lumberyards[2297]}));
acre acre_45_48 (.clk(clk), .en(en), .top_left({trees[2247], lumberyards[2247]}), .top({trees[2248], lumberyards[2248]}), .top_right({trees[2249], lumberyards[2249]}), .left({trees[2297], lumberyards[2297]}), .right({trees[2299], lumberyards[2299]}), .bottom_left({trees[2347], lumberyards[2347]}), .bottom({trees[2348], lumberyards[2348]}), .bottom_right({trees[2349], lumberyards[2349]}), .init(2'b00), .state({trees[2298], lumberyards[2298]}));
acre acre_45_49 (.clk(clk), .en(en), .top_left({trees[2248], lumberyards[2248]}), .top({trees[2249], lumberyards[2249]}), .top_right(2'b0), .left({trees[2298], lumberyards[2298]}), .right(2'b0), .bottom_left({trees[2348], lumberyards[2348]}), .bottom({trees[2349], lumberyards[2349]}), .bottom_right(2'b0), .init(2'b00), .state({trees[2299], lumberyards[2299]}));
acre acre_46_0 (.clk(clk), .en(en), .top_left(2'b0), .top({trees[2250], lumberyards[2250]}), .top_right({trees[2251], lumberyards[2251]}), .left(2'b0), .right({trees[2301], lumberyards[2301]}), .bottom_left(2'b0), .bottom({trees[2350], lumberyards[2350]}), .bottom_right({trees[2351], lumberyards[2351]}), .init(2'b10), .state({trees[2300], lumberyards[2300]}));
acre acre_46_1 (.clk(clk), .en(en), .top_left({trees[2250], lumberyards[2250]}), .top({trees[2251], lumberyards[2251]}), .top_right({trees[2252], lumberyards[2252]}), .left({trees[2300], lumberyards[2300]}), .right({trees[2302], lumberyards[2302]}), .bottom_left({trees[2350], lumberyards[2350]}), .bottom({trees[2351], lumberyards[2351]}), .bottom_right({trees[2352], lumberyards[2352]}), .init(2'b10), .state({trees[2301], lumberyards[2301]}));
acre acre_46_2 (.clk(clk), .en(en), .top_left({trees[2251], lumberyards[2251]}), .top({trees[2252], lumberyards[2252]}), .top_right({trees[2253], lumberyards[2253]}), .left({trees[2301], lumberyards[2301]}), .right({trees[2303], lumberyards[2303]}), .bottom_left({trees[2351], lumberyards[2351]}), .bottom({trees[2352], lumberyards[2352]}), .bottom_right({trees[2353], lumberyards[2353]}), .init(2'b00), .state({trees[2302], lumberyards[2302]}));
acre acre_46_3 (.clk(clk), .en(en), .top_left({trees[2252], lumberyards[2252]}), .top({trees[2253], lumberyards[2253]}), .top_right({trees[2254], lumberyards[2254]}), .left({trees[2302], lumberyards[2302]}), .right({trees[2304], lumberyards[2304]}), .bottom_left({trees[2352], lumberyards[2352]}), .bottom({trees[2353], lumberyards[2353]}), .bottom_right({trees[2354], lumberyards[2354]}), .init(2'b00), .state({trees[2303], lumberyards[2303]}));
acre acre_46_4 (.clk(clk), .en(en), .top_left({trees[2253], lumberyards[2253]}), .top({trees[2254], lumberyards[2254]}), .top_right({trees[2255], lumberyards[2255]}), .left({trees[2303], lumberyards[2303]}), .right({trees[2305], lumberyards[2305]}), .bottom_left({trees[2353], lumberyards[2353]}), .bottom({trees[2354], lumberyards[2354]}), .bottom_right({trees[2355], lumberyards[2355]}), .init(2'b01), .state({trees[2304], lumberyards[2304]}));
acre acre_46_5 (.clk(clk), .en(en), .top_left({trees[2254], lumberyards[2254]}), .top({trees[2255], lumberyards[2255]}), .top_right({trees[2256], lumberyards[2256]}), .left({trees[2304], lumberyards[2304]}), .right({trees[2306], lumberyards[2306]}), .bottom_left({trees[2354], lumberyards[2354]}), .bottom({trees[2355], lumberyards[2355]}), .bottom_right({trees[2356], lumberyards[2356]}), .init(2'b00), .state({trees[2305], lumberyards[2305]}));
acre acre_46_6 (.clk(clk), .en(en), .top_left({trees[2255], lumberyards[2255]}), .top({trees[2256], lumberyards[2256]}), .top_right({trees[2257], lumberyards[2257]}), .left({trees[2305], lumberyards[2305]}), .right({trees[2307], lumberyards[2307]}), .bottom_left({trees[2355], lumberyards[2355]}), .bottom({trees[2356], lumberyards[2356]}), .bottom_right({trees[2357], lumberyards[2357]}), .init(2'b01), .state({trees[2306], lumberyards[2306]}));
acre acre_46_7 (.clk(clk), .en(en), .top_left({trees[2256], lumberyards[2256]}), .top({trees[2257], lumberyards[2257]}), .top_right({trees[2258], lumberyards[2258]}), .left({trees[2306], lumberyards[2306]}), .right({trees[2308], lumberyards[2308]}), .bottom_left({trees[2356], lumberyards[2356]}), .bottom({trees[2357], lumberyards[2357]}), .bottom_right({trees[2358], lumberyards[2358]}), .init(2'b10), .state({trees[2307], lumberyards[2307]}));
acre acre_46_8 (.clk(clk), .en(en), .top_left({trees[2257], lumberyards[2257]}), .top({trees[2258], lumberyards[2258]}), .top_right({trees[2259], lumberyards[2259]}), .left({trees[2307], lumberyards[2307]}), .right({trees[2309], lumberyards[2309]}), .bottom_left({trees[2357], lumberyards[2357]}), .bottom({trees[2358], lumberyards[2358]}), .bottom_right({trees[2359], lumberyards[2359]}), .init(2'b00), .state({trees[2308], lumberyards[2308]}));
acre acre_46_9 (.clk(clk), .en(en), .top_left({trees[2258], lumberyards[2258]}), .top({trees[2259], lumberyards[2259]}), .top_right({trees[2260], lumberyards[2260]}), .left({trees[2308], lumberyards[2308]}), .right({trees[2310], lumberyards[2310]}), .bottom_left({trees[2358], lumberyards[2358]}), .bottom({trees[2359], lumberyards[2359]}), .bottom_right({trees[2360], lumberyards[2360]}), .init(2'b00), .state({trees[2309], lumberyards[2309]}));
acre acre_46_10 (.clk(clk), .en(en), .top_left({trees[2259], lumberyards[2259]}), .top({trees[2260], lumberyards[2260]}), .top_right({trees[2261], lumberyards[2261]}), .left({trees[2309], lumberyards[2309]}), .right({trees[2311], lumberyards[2311]}), .bottom_left({trees[2359], lumberyards[2359]}), .bottom({trees[2360], lumberyards[2360]}), .bottom_right({trees[2361], lumberyards[2361]}), .init(2'b10), .state({trees[2310], lumberyards[2310]}));
acre acre_46_11 (.clk(clk), .en(en), .top_left({trees[2260], lumberyards[2260]}), .top({trees[2261], lumberyards[2261]}), .top_right({trees[2262], lumberyards[2262]}), .left({trees[2310], lumberyards[2310]}), .right({trees[2312], lumberyards[2312]}), .bottom_left({trees[2360], lumberyards[2360]}), .bottom({trees[2361], lumberyards[2361]}), .bottom_right({trees[2362], lumberyards[2362]}), .init(2'b00), .state({trees[2311], lumberyards[2311]}));
acre acre_46_12 (.clk(clk), .en(en), .top_left({trees[2261], lumberyards[2261]}), .top({trees[2262], lumberyards[2262]}), .top_right({trees[2263], lumberyards[2263]}), .left({trees[2311], lumberyards[2311]}), .right({trees[2313], lumberyards[2313]}), .bottom_left({trees[2361], lumberyards[2361]}), .bottom({trees[2362], lumberyards[2362]}), .bottom_right({trees[2363], lumberyards[2363]}), .init(2'b10), .state({trees[2312], lumberyards[2312]}));
acre acre_46_13 (.clk(clk), .en(en), .top_left({trees[2262], lumberyards[2262]}), .top({trees[2263], lumberyards[2263]}), .top_right({trees[2264], lumberyards[2264]}), .left({trees[2312], lumberyards[2312]}), .right({trees[2314], lumberyards[2314]}), .bottom_left({trees[2362], lumberyards[2362]}), .bottom({trees[2363], lumberyards[2363]}), .bottom_right({trees[2364], lumberyards[2364]}), .init(2'b01), .state({trees[2313], lumberyards[2313]}));
acre acre_46_14 (.clk(clk), .en(en), .top_left({trees[2263], lumberyards[2263]}), .top({trees[2264], lumberyards[2264]}), .top_right({trees[2265], lumberyards[2265]}), .left({trees[2313], lumberyards[2313]}), .right({trees[2315], lumberyards[2315]}), .bottom_left({trees[2363], lumberyards[2363]}), .bottom({trees[2364], lumberyards[2364]}), .bottom_right({trees[2365], lumberyards[2365]}), .init(2'b00), .state({trees[2314], lumberyards[2314]}));
acre acre_46_15 (.clk(clk), .en(en), .top_left({trees[2264], lumberyards[2264]}), .top({trees[2265], lumberyards[2265]}), .top_right({trees[2266], lumberyards[2266]}), .left({trees[2314], lumberyards[2314]}), .right({trees[2316], lumberyards[2316]}), .bottom_left({trees[2364], lumberyards[2364]}), .bottom({trees[2365], lumberyards[2365]}), .bottom_right({trees[2366], lumberyards[2366]}), .init(2'b00), .state({trees[2315], lumberyards[2315]}));
acre acre_46_16 (.clk(clk), .en(en), .top_left({trees[2265], lumberyards[2265]}), .top({trees[2266], lumberyards[2266]}), .top_right({trees[2267], lumberyards[2267]}), .left({trees[2315], lumberyards[2315]}), .right({trees[2317], lumberyards[2317]}), .bottom_left({trees[2365], lumberyards[2365]}), .bottom({trees[2366], lumberyards[2366]}), .bottom_right({trees[2367], lumberyards[2367]}), .init(2'b10), .state({trees[2316], lumberyards[2316]}));
acre acre_46_17 (.clk(clk), .en(en), .top_left({trees[2266], lumberyards[2266]}), .top({trees[2267], lumberyards[2267]}), .top_right({trees[2268], lumberyards[2268]}), .left({trees[2316], lumberyards[2316]}), .right({trees[2318], lumberyards[2318]}), .bottom_left({trees[2366], lumberyards[2366]}), .bottom({trees[2367], lumberyards[2367]}), .bottom_right({trees[2368], lumberyards[2368]}), .init(2'b00), .state({trees[2317], lumberyards[2317]}));
acre acre_46_18 (.clk(clk), .en(en), .top_left({trees[2267], lumberyards[2267]}), .top({trees[2268], lumberyards[2268]}), .top_right({trees[2269], lumberyards[2269]}), .left({trees[2317], lumberyards[2317]}), .right({trees[2319], lumberyards[2319]}), .bottom_left({trees[2367], lumberyards[2367]}), .bottom({trees[2368], lumberyards[2368]}), .bottom_right({trees[2369], lumberyards[2369]}), .init(2'b00), .state({trees[2318], lumberyards[2318]}));
acre acre_46_19 (.clk(clk), .en(en), .top_left({trees[2268], lumberyards[2268]}), .top({trees[2269], lumberyards[2269]}), .top_right({trees[2270], lumberyards[2270]}), .left({trees[2318], lumberyards[2318]}), .right({trees[2320], lumberyards[2320]}), .bottom_left({trees[2368], lumberyards[2368]}), .bottom({trees[2369], lumberyards[2369]}), .bottom_right({trees[2370], lumberyards[2370]}), .init(2'b00), .state({trees[2319], lumberyards[2319]}));
acre acre_46_20 (.clk(clk), .en(en), .top_left({trees[2269], lumberyards[2269]}), .top({trees[2270], lumberyards[2270]}), .top_right({trees[2271], lumberyards[2271]}), .left({trees[2319], lumberyards[2319]}), .right({trees[2321], lumberyards[2321]}), .bottom_left({trees[2369], lumberyards[2369]}), .bottom({trees[2370], lumberyards[2370]}), .bottom_right({trees[2371], lumberyards[2371]}), .init(2'b01), .state({trees[2320], lumberyards[2320]}));
acre acre_46_21 (.clk(clk), .en(en), .top_left({trees[2270], lumberyards[2270]}), .top({trees[2271], lumberyards[2271]}), .top_right({trees[2272], lumberyards[2272]}), .left({trees[2320], lumberyards[2320]}), .right({trees[2322], lumberyards[2322]}), .bottom_left({trees[2370], lumberyards[2370]}), .bottom({trees[2371], lumberyards[2371]}), .bottom_right({trees[2372], lumberyards[2372]}), .init(2'b01), .state({trees[2321], lumberyards[2321]}));
acre acre_46_22 (.clk(clk), .en(en), .top_left({trees[2271], lumberyards[2271]}), .top({trees[2272], lumberyards[2272]}), .top_right({trees[2273], lumberyards[2273]}), .left({trees[2321], lumberyards[2321]}), .right({trees[2323], lumberyards[2323]}), .bottom_left({trees[2371], lumberyards[2371]}), .bottom({trees[2372], lumberyards[2372]}), .bottom_right({trees[2373], lumberyards[2373]}), .init(2'b00), .state({trees[2322], lumberyards[2322]}));
acre acre_46_23 (.clk(clk), .en(en), .top_left({trees[2272], lumberyards[2272]}), .top({trees[2273], lumberyards[2273]}), .top_right({trees[2274], lumberyards[2274]}), .left({trees[2322], lumberyards[2322]}), .right({trees[2324], lumberyards[2324]}), .bottom_left({trees[2372], lumberyards[2372]}), .bottom({trees[2373], lumberyards[2373]}), .bottom_right({trees[2374], lumberyards[2374]}), .init(2'b00), .state({trees[2323], lumberyards[2323]}));
acre acre_46_24 (.clk(clk), .en(en), .top_left({trees[2273], lumberyards[2273]}), .top({trees[2274], lumberyards[2274]}), .top_right({trees[2275], lumberyards[2275]}), .left({trees[2323], lumberyards[2323]}), .right({trees[2325], lumberyards[2325]}), .bottom_left({trees[2373], lumberyards[2373]}), .bottom({trees[2374], lumberyards[2374]}), .bottom_right({trees[2375], lumberyards[2375]}), .init(2'b00), .state({trees[2324], lumberyards[2324]}));
acre acre_46_25 (.clk(clk), .en(en), .top_left({trees[2274], lumberyards[2274]}), .top({trees[2275], lumberyards[2275]}), .top_right({trees[2276], lumberyards[2276]}), .left({trees[2324], lumberyards[2324]}), .right({trees[2326], lumberyards[2326]}), .bottom_left({trees[2374], lumberyards[2374]}), .bottom({trees[2375], lumberyards[2375]}), .bottom_right({trees[2376], lumberyards[2376]}), .init(2'b00), .state({trees[2325], lumberyards[2325]}));
acre acre_46_26 (.clk(clk), .en(en), .top_left({trees[2275], lumberyards[2275]}), .top({trees[2276], lumberyards[2276]}), .top_right({trees[2277], lumberyards[2277]}), .left({trees[2325], lumberyards[2325]}), .right({trees[2327], lumberyards[2327]}), .bottom_left({trees[2375], lumberyards[2375]}), .bottom({trees[2376], lumberyards[2376]}), .bottom_right({trees[2377], lumberyards[2377]}), .init(2'b00), .state({trees[2326], lumberyards[2326]}));
acre acre_46_27 (.clk(clk), .en(en), .top_left({trees[2276], lumberyards[2276]}), .top({trees[2277], lumberyards[2277]}), .top_right({trees[2278], lumberyards[2278]}), .left({trees[2326], lumberyards[2326]}), .right({trees[2328], lumberyards[2328]}), .bottom_left({trees[2376], lumberyards[2376]}), .bottom({trees[2377], lumberyards[2377]}), .bottom_right({trees[2378], lumberyards[2378]}), .init(2'b00), .state({trees[2327], lumberyards[2327]}));
acre acre_46_28 (.clk(clk), .en(en), .top_left({trees[2277], lumberyards[2277]}), .top({trees[2278], lumberyards[2278]}), .top_right({trees[2279], lumberyards[2279]}), .left({trees[2327], lumberyards[2327]}), .right({trees[2329], lumberyards[2329]}), .bottom_left({trees[2377], lumberyards[2377]}), .bottom({trees[2378], lumberyards[2378]}), .bottom_right({trees[2379], lumberyards[2379]}), .init(2'b00), .state({trees[2328], lumberyards[2328]}));
acre acre_46_29 (.clk(clk), .en(en), .top_left({trees[2278], lumberyards[2278]}), .top({trees[2279], lumberyards[2279]}), .top_right({trees[2280], lumberyards[2280]}), .left({trees[2328], lumberyards[2328]}), .right({trees[2330], lumberyards[2330]}), .bottom_left({trees[2378], lumberyards[2378]}), .bottom({trees[2379], lumberyards[2379]}), .bottom_right({trees[2380], lumberyards[2380]}), .init(2'b00), .state({trees[2329], lumberyards[2329]}));
acre acre_46_30 (.clk(clk), .en(en), .top_left({trees[2279], lumberyards[2279]}), .top({trees[2280], lumberyards[2280]}), .top_right({trees[2281], lumberyards[2281]}), .left({trees[2329], lumberyards[2329]}), .right({trees[2331], lumberyards[2331]}), .bottom_left({trees[2379], lumberyards[2379]}), .bottom({trees[2380], lumberyards[2380]}), .bottom_right({trees[2381], lumberyards[2381]}), .init(2'b00), .state({trees[2330], lumberyards[2330]}));
acre acre_46_31 (.clk(clk), .en(en), .top_left({trees[2280], lumberyards[2280]}), .top({trees[2281], lumberyards[2281]}), .top_right({trees[2282], lumberyards[2282]}), .left({trees[2330], lumberyards[2330]}), .right({trees[2332], lumberyards[2332]}), .bottom_left({trees[2380], lumberyards[2380]}), .bottom({trees[2381], lumberyards[2381]}), .bottom_right({trees[2382], lumberyards[2382]}), .init(2'b00), .state({trees[2331], lumberyards[2331]}));
acre acre_46_32 (.clk(clk), .en(en), .top_left({trees[2281], lumberyards[2281]}), .top({trees[2282], lumberyards[2282]}), .top_right({trees[2283], lumberyards[2283]}), .left({trees[2331], lumberyards[2331]}), .right({trees[2333], lumberyards[2333]}), .bottom_left({trees[2381], lumberyards[2381]}), .bottom({trees[2382], lumberyards[2382]}), .bottom_right({trees[2383], lumberyards[2383]}), .init(2'b00), .state({trees[2332], lumberyards[2332]}));
acre acre_46_33 (.clk(clk), .en(en), .top_left({trees[2282], lumberyards[2282]}), .top({trees[2283], lumberyards[2283]}), .top_right({trees[2284], lumberyards[2284]}), .left({trees[2332], lumberyards[2332]}), .right({trees[2334], lumberyards[2334]}), .bottom_left({trees[2382], lumberyards[2382]}), .bottom({trees[2383], lumberyards[2383]}), .bottom_right({trees[2384], lumberyards[2384]}), .init(2'b01), .state({trees[2333], lumberyards[2333]}));
acre acre_46_34 (.clk(clk), .en(en), .top_left({trees[2283], lumberyards[2283]}), .top({trees[2284], lumberyards[2284]}), .top_right({trees[2285], lumberyards[2285]}), .left({trees[2333], lumberyards[2333]}), .right({trees[2335], lumberyards[2335]}), .bottom_left({trees[2383], lumberyards[2383]}), .bottom({trees[2384], lumberyards[2384]}), .bottom_right({trees[2385], lumberyards[2385]}), .init(2'b00), .state({trees[2334], lumberyards[2334]}));
acre acre_46_35 (.clk(clk), .en(en), .top_left({trees[2284], lumberyards[2284]}), .top({trees[2285], lumberyards[2285]}), .top_right({trees[2286], lumberyards[2286]}), .left({trees[2334], lumberyards[2334]}), .right({trees[2336], lumberyards[2336]}), .bottom_left({trees[2384], lumberyards[2384]}), .bottom({trees[2385], lumberyards[2385]}), .bottom_right({trees[2386], lumberyards[2386]}), .init(2'b10), .state({trees[2335], lumberyards[2335]}));
acre acre_46_36 (.clk(clk), .en(en), .top_left({trees[2285], lumberyards[2285]}), .top({trees[2286], lumberyards[2286]}), .top_right({trees[2287], lumberyards[2287]}), .left({trees[2335], lumberyards[2335]}), .right({trees[2337], lumberyards[2337]}), .bottom_left({trees[2385], lumberyards[2385]}), .bottom({trees[2386], lumberyards[2386]}), .bottom_right({trees[2387], lumberyards[2387]}), .init(2'b10), .state({trees[2336], lumberyards[2336]}));
acre acre_46_37 (.clk(clk), .en(en), .top_left({trees[2286], lumberyards[2286]}), .top({trees[2287], lumberyards[2287]}), .top_right({trees[2288], lumberyards[2288]}), .left({trees[2336], lumberyards[2336]}), .right({trees[2338], lumberyards[2338]}), .bottom_left({trees[2386], lumberyards[2386]}), .bottom({trees[2387], lumberyards[2387]}), .bottom_right({trees[2388], lumberyards[2388]}), .init(2'b00), .state({trees[2337], lumberyards[2337]}));
acre acre_46_38 (.clk(clk), .en(en), .top_left({trees[2287], lumberyards[2287]}), .top({trees[2288], lumberyards[2288]}), .top_right({trees[2289], lumberyards[2289]}), .left({trees[2337], lumberyards[2337]}), .right({trees[2339], lumberyards[2339]}), .bottom_left({trees[2387], lumberyards[2387]}), .bottom({trees[2388], lumberyards[2388]}), .bottom_right({trees[2389], lumberyards[2389]}), .init(2'b10), .state({trees[2338], lumberyards[2338]}));
acre acre_46_39 (.clk(clk), .en(en), .top_left({trees[2288], lumberyards[2288]}), .top({trees[2289], lumberyards[2289]}), .top_right({trees[2290], lumberyards[2290]}), .left({trees[2338], lumberyards[2338]}), .right({trees[2340], lumberyards[2340]}), .bottom_left({trees[2388], lumberyards[2388]}), .bottom({trees[2389], lumberyards[2389]}), .bottom_right({trees[2390], lumberyards[2390]}), .init(2'b00), .state({trees[2339], lumberyards[2339]}));
acre acre_46_40 (.clk(clk), .en(en), .top_left({trees[2289], lumberyards[2289]}), .top({trees[2290], lumberyards[2290]}), .top_right({trees[2291], lumberyards[2291]}), .left({trees[2339], lumberyards[2339]}), .right({trees[2341], lumberyards[2341]}), .bottom_left({trees[2389], lumberyards[2389]}), .bottom({trees[2390], lumberyards[2390]}), .bottom_right({trees[2391], lumberyards[2391]}), .init(2'b00), .state({trees[2340], lumberyards[2340]}));
acre acre_46_41 (.clk(clk), .en(en), .top_left({trees[2290], lumberyards[2290]}), .top({trees[2291], lumberyards[2291]}), .top_right({trees[2292], lumberyards[2292]}), .left({trees[2340], lumberyards[2340]}), .right({trees[2342], lumberyards[2342]}), .bottom_left({trees[2390], lumberyards[2390]}), .bottom({trees[2391], lumberyards[2391]}), .bottom_right({trees[2392], lumberyards[2392]}), .init(2'b01), .state({trees[2341], lumberyards[2341]}));
acre acre_46_42 (.clk(clk), .en(en), .top_left({trees[2291], lumberyards[2291]}), .top({trees[2292], lumberyards[2292]}), .top_right({trees[2293], lumberyards[2293]}), .left({trees[2341], lumberyards[2341]}), .right({trees[2343], lumberyards[2343]}), .bottom_left({trees[2391], lumberyards[2391]}), .bottom({trees[2392], lumberyards[2392]}), .bottom_right({trees[2393], lumberyards[2393]}), .init(2'b01), .state({trees[2342], lumberyards[2342]}));
acre acre_46_43 (.clk(clk), .en(en), .top_left({trees[2292], lumberyards[2292]}), .top({trees[2293], lumberyards[2293]}), .top_right({trees[2294], lumberyards[2294]}), .left({trees[2342], lumberyards[2342]}), .right({trees[2344], lumberyards[2344]}), .bottom_left({trees[2392], lumberyards[2392]}), .bottom({trees[2393], lumberyards[2393]}), .bottom_right({trees[2394], lumberyards[2394]}), .init(2'b00), .state({trees[2343], lumberyards[2343]}));
acre acre_46_44 (.clk(clk), .en(en), .top_left({trees[2293], lumberyards[2293]}), .top({trees[2294], lumberyards[2294]}), .top_right({trees[2295], lumberyards[2295]}), .left({trees[2343], lumberyards[2343]}), .right({trees[2345], lumberyards[2345]}), .bottom_left({trees[2393], lumberyards[2393]}), .bottom({trees[2394], lumberyards[2394]}), .bottom_right({trees[2395], lumberyards[2395]}), .init(2'b00), .state({trees[2344], lumberyards[2344]}));
acre acre_46_45 (.clk(clk), .en(en), .top_left({trees[2294], lumberyards[2294]}), .top({trees[2295], lumberyards[2295]}), .top_right({trees[2296], lumberyards[2296]}), .left({trees[2344], lumberyards[2344]}), .right({trees[2346], lumberyards[2346]}), .bottom_left({trees[2394], lumberyards[2394]}), .bottom({trees[2395], lumberyards[2395]}), .bottom_right({trees[2396], lumberyards[2396]}), .init(2'b01), .state({trees[2345], lumberyards[2345]}));
acre acre_46_46 (.clk(clk), .en(en), .top_left({trees[2295], lumberyards[2295]}), .top({trees[2296], lumberyards[2296]}), .top_right({trees[2297], lumberyards[2297]}), .left({trees[2345], lumberyards[2345]}), .right({trees[2347], lumberyards[2347]}), .bottom_left({trees[2395], lumberyards[2395]}), .bottom({trees[2396], lumberyards[2396]}), .bottom_right({trees[2397], lumberyards[2397]}), .init(2'b00), .state({trees[2346], lumberyards[2346]}));
acre acre_46_47 (.clk(clk), .en(en), .top_left({trees[2296], lumberyards[2296]}), .top({trees[2297], lumberyards[2297]}), .top_right({trees[2298], lumberyards[2298]}), .left({trees[2346], lumberyards[2346]}), .right({trees[2348], lumberyards[2348]}), .bottom_left({trees[2396], lumberyards[2396]}), .bottom({trees[2397], lumberyards[2397]}), .bottom_right({trees[2398], lumberyards[2398]}), .init(2'b10), .state({trees[2347], lumberyards[2347]}));
acre acre_46_48 (.clk(clk), .en(en), .top_left({trees[2297], lumberyards[2297]}), .top({trees[2298], lumberyards[2298]}), .top_right({trees[2299], lumberyards[2299]}), .left({trees[2347], lumberyards[2347]}), .right({trees[2349], lumberyards[2349]}), .bottom_left({trees[2397], lumberyards[2397]}), .bottom({trees[2398], lumberyards[2398]}), .bottom_right({trees[2399], lumberyards[2399]}), .init(2'b00), .state({trees[2348], lumberyards[2348]}));
acre acre_46_49 (.clk(clk), .en(en), .top_left({trees[2298], lumberyards[2298]}), .top({trees[2299], lumberyards[2299]}), .top_right(2'b0), .left({trees[2348], lumberyards[2348]}), .right(2'b0), .bottom_left({trees[2398], lumberyards[2398]}), .bottom({trees[2399], lumberyards[2399]}), .bottom_right(2'b0), .init(2'b00), .state({trees[2349], lumberyards[2349]}));
acre acre_47_0 (.clk(clk), .en(en), .top_left(2'b0), .top({trees[2300], lumberyards[2300]}), .top_right({trees[2301], lumberyards[2301]}), .left(2'b0), .right({trees[2351], lumberyards[2351]}), .bottom_left(2'b0), .bottom({trees[2400], lumberyards[2400]}), .bottom_right({trees[2401], lumberyards[2401]}), .init(2'b00), .state({trees[2350], lumberyards[2350]}));
acre acre_47_1 (.clk(clk), .en(en), .top_left({trees[2300], lumberyards[2300]}), .top({trees[2301], lumberyards[2301]}), .top_right({trees[2302], lumberyards[2302]}), .left({trees[2350], lumberyards[2350]}), .right({trees[2352], lumberyards[2352]}), .bottom_left({trees[2400], lumberyards[2400]}), .bottom({trees[2401], lumberyards[2401]}), .bottom_right({trees[2402], lumberyards[2402]}), .init(2'b00), .state({trees[2351], lumberyards[2351]}));
acre acre_47_2 (.clk(clk), .en(en), .top_left({trees[2301], lumberyards[2301]}), .top({trees[2302], lumberyards[2302]}), .top_right({trees[2303], lumberyards[2303]}), .left({trees[2351], lumberyards[2351]}), .right({trees[2353], lumberyards[2353]}), .bottom_left({trees[2401], lumberyards[2401]}), .bottom({trees[2402], lumberyards[2402]}), .bottom_right({trees[2403], lumberyards[2403]}), .init(2'b00), .state({trees[2352], lumberyards[2352]}));
acre acre_47_3 (.clk(clk), .en(en), .top_left({trees[2302], lumberyards[2302]}), .top({trees[2303], lumberyards[2303]}), .top_right({trees[2304], lumberyards[2304]}), .left({trees[2352], lumberyards[2352]}), .right({trees[2354], lumberyards[2354]}), .bottom_left({trees[2402], lumberyards[2402]}), .bottom({trees[2403], lumberyards[2403]}), .bottom_right({trees[2404], lumberyards[2404]}), .init(2'b00), .state({trees[2353], lumberyards[2353]}));
acre acre_47_4 (.clk(clk), .en(en), .top_left({trees[2303], lumberyards[2303]}), .top({trees[2304], lumberyards[2304]}), .top_right({trees[2305], lumberyards[2305]}), .left({trees[2353], lumberyards[2353]}), .right({trees[2355], lumberyards[2355]}), .bottom_left({trees[2403], lumberyards[2403]}), .bottom({trees[2404], lumberyards[2404]}), .bottom_right({trees[2405], lumberyards[2405]}), .init(2'b00), .state({trees[2354], lumberyards[2354]}));
acre acre_47_5 (.clk(clk), .en(en), .top_left({trees[2304], lumberyards[2304]}), .top({trees[2305], lumberyards[2305]}), .top_right({trees[2306], lumberyards[2306]}), .left({trees[2354], lumberyards[2354]}), .right({trees[2356], lumberyards[2356]}), .bottom_left({trees[2404], lumberyards[2404]}), .bottom({trees[2405], lumberyards[2405]}), .bottom_right({trees[2406], lumberyards[2406]}), .init(2'b00), .state({trees[2355], lumberyards[2355]}));
acre acre_47_6 (.clk(clk), .en(en), .top_left({trees[2305], lumberyards[2305]}), .top({trees[2306], lumberyards[2306]}), .top_right({trees[2307], lumberyards[2307]}), .left({trees[2355], lumberyards[2355]}), .right({trees[2357], lumberyards[2357]}), .bottom_left({trees[2405], lumberyards[2405]}), .bottom({trees[2406], lumberyards[2406]}), .bottom_right({trees[2407], lumberyards[2407]}), .init(2'b00), .state({trees[2356], lumberyards[2356]}));
acre acre_47_7 (.clk(clk), .en(en), .top_left({trees[2306], lumberyards[2306]}), .top({trees[2307], lumberyards[2307]}), .top_right({trees[2308], lumberyards[2308]}), .left({trees[2356], lumberyards[2356]}), .right({trees[2358], lumberyards[2358]}), .bottom_left({trees[2406], lumberyards[2406]}), .bottom({trees[2407], lumberyards[2407]}), .bottom_right({trees[2408], lumberyards[2408]}), .init(2'b10), .state({trees[2357], lumberyards[2357]}));
acre acre_47_8 (.clk(clk), .en(en), .top_left({trees[2307], lumberyards[2307]}), .top({trees[2308], lumberyards[2308]}), .top_right({trees[2309], lumberyards[2309]}), .left({trees[2357], lumberyards[2357]}), .right({trees[2359], lumberyards[2359]}), .bottom_left({trees[2407], lumberyards[2407]}), .bottom({trees[2408], lumberyards[2408]}), .bottom_right({trees[2409], lumberyards[2409]}), .init(2'b00), .state({trees[2358], lumberyards[2358]}));
acre acre_47_9 (.clk(clk), .en(en), .top_left({trees[2308], lumberyards[2308]}), .top({trees[2309], lumberyards[2309]}), .top_right({trees[2310], lumberyards[2310]}), .left({trees[2358], lumberyards[2358]}), .right({trees[2360], lumberyards[2360]}), .bottom_left({trees[2408], lumberyards[2408]}), .bottom({trees[2409], lumberyards[2409]}), .bottom_right({trees[2410], lumberyards[2410]}), .init(2'b10), .state({trees[2359], lumberyards[2359]}));
acre acre_47_10 (.clk(clk), .en(en), .top_left({trees[2309], lumberyards[2309]}), .top({trees[2310], lumberyards[2310]}), .top_right({trees[2311], lumberyards[2311]}), .left({trees[2359], lumberyards[2359]}), .right({trees[2361], lumberyards[2361]}), .bottom_left({trees[2409], lumberyards[2409]}), .bottom({trees[2410], lumberyards[2410]}), .bottom_right({trees[2411], lumberyards[2411]}), .init(2'b00), .state({trees[2360], lumberyards[2360]}));
acre acre_47_11 (.clk(clk), .en(en), .top_left({trees[2310], lumberyards[2310]}), .top({trees[2311], lumberyards[2311]}), .top_right({trees[2312], lumberyards[2312]}), .left({trees[2360], lumberyards[2360]}), .right({trees[2362], lumberyards[2362]}), .bottom_left({trees[2410], lumberyards[2410]}), .bottom({trees[2411], lumberyards[2411]}), .bottom_right({trees[2412], lumberyards[2412]}), .init(2'b10), .state({trees[2361], lumberyards[2361]}));
acre acre_47_12 (.clk(clk), .en(en), .top_left({trees[2311], lumberyards[2311]}), .top({trees[2312], lumberyards[2312]}), .top_right({trees[2313], lumberyards[2313]}), .left({trees[2361], lumberyards[2361]}), .right({trees[2363], lumberyards[2363]}), .bottom_left({trees[2411], lumberyards[2411]}), .bottom({trees[2412], lumberyards[2412]}), .bottom_right({trees[2413], lumberyards[2413]}), .init(2'b00), .state({trees[2362], lumberyards[2362]}));
acre acre_47_13 (.clk(clk), .en(en), .top_left({trees[2312], lumberyards[2312]}), .top({trees[2313], lumberyards[2313]}), .top_right({trees[2314], lumberyards[2314]}), .left({trees[2362], lumberyards[2362]}), .right({trees[2364], lumberyards[2364]}), .bottom_left({trees[2412], lumberyards[2412]}), .bottom({trees[2413], lumberyards[2413]}), .bottom_right({trees[2414], lumberyards[2414]}), .init(2'b00), .state({trees[2363], lumberyards[2363]}));
acre acre_47_14 (.clk(clk), .en(en), .top_left({trees[2313], lumberyards[2313]}), .top({trees[2314], lumberyards[2314]}), .top_right({trees[2315], lumberyards[2315]}), .left({trees[2363], lumberyards[2363]}), .right({trees[2365], lumberyards[2365]}), .bottom_left({trees[2413], lumberyards[2413]}), .bottom({trees[2414], lumberyards[2414]}), .bottom_right({trees[2415], lumberyards[2415]}), .init(2'b00), .state({trees[2364], lumberyards[2364]}));
acre acre_47_15 (.clk(clk), .en(en), .top_left({trees[2314], lumberyards[2314]}), .top({trees[2315], lumberyards[2315]}), .top_right({trees[2316], lumberyards[2316]}), .left({trees[2364], lumberyards[2364]}), .right({trees[2366], lumberyards[2366]}), .bottom_left({trees[2414], lumberyards[2414]}), .bottom({trees[2415], lumberyards[2415]}), .bottom_right({trees[2416], lumberyards[2416]}), .init(2'b10), .state({trees[2365], lumberyards[2365]}));
acre acre_47_16 (.clk(clk), .en(en), .top_left({trees[2315], lumberyards[2315]}), .top({trees[2316], lumberyards[2316]}), .top_right({trees[2317], lumberyards[2317]}), .left({trees[2365], lumberyards[2365]}), .right({trees[2367], lumberyards[2367]}), .bottom_left({trees[2415], lumberyards[2415]}), .bottom({trees[2416], lumberyards[2416]}), .bottom_right({trees[2417], lumberyards[2417]}), .init(2'b00), .state({trees[2366], lumberyards[2366]}));
acre acre_47_17 (.clk(clk), .en(en), .top_left({trees[2316], lumberyards[2316]}), .top({trees[2317], lumberyards[2317]}), .top_right({trees[2318], lumberyards[2318]}), .left({trees[2366], lumberyards[2366]}), .right({trees[2368], lumberyards[2368]}), .bottom_left({trees[2416], lumberyards[2416]}), .bottom({trees[2417], lumberyards[2417]}), .bottom_right({trees[2418], lumberyards[2418]}), .init(2'b00), .state({trees[2367], lumberyards[2367]}));
acre acre_47_18 (.clk(clk), .en(en), .top_left({trees[2317], lumberyards[2317]}), .top({trees[2318], lumberyards[2318]}), .top_right({trees[2319], lumberyards[2319]}), .left({trees[2367], lumberyards[2367]}), .right({trees[2369], lumberyards[2369]}), .bottom_left({trees[2417], lumberyards[2417]}), .bottom({trees[2418], lumberyards[2418]}), .bottom_right({trees[2419], lumberyards[2419]}), .init(2'b00), .state({trees[2368], lumberyards[2368]}));
acre acre_47_19 (.clk(clk), .en(en), .top_left({trees[2318], lumberyards[2318]}), .top({trees[2319], lumberyards[2319]}), .top_right({trees[2320], lumberyards[2320]}), .left({trees[2368], lumberyards[2368]}), .right({trees[2370], lumberyards[2370]}), .bottom_left({trees[2418], lumberyards[2418]}), .bottom({trees[2419], lumberyards[2419]}), .bottom_right({trees[2420], lumberyards[2420]}), .init(2'b01), .state({trees[2369], lumberyards[2369]}));
acre acre_47_20 (.clk(clk), .en(en), .top_left({trees[2319], lumberyards[2319]}), .top({trees[2320], lumberyards[2320]}), .top_right({trees[2321], lumberyards[2321]}), .left({trees[2369], lumberyards[2369]}), .right({trees[2371], lumberyards[2371]}), .bottom_left({trees[2419], lumberyards[2419]}), .bottom({trees[2420], lumberyards[2420]}), .bottom_right({trees[2421], lumberyards[2421]}), .init(2'b00), .state({trees[2370], lumberyards[2370]}));
acre acre_47_21 (.clk(clk), .en(en), .top_left({trees[2320], lumberyards[2320]}), .top({trees[2321], lumberyards[2321]}), .top_right({trees[2322], lumberyards[2322]}), .left({trees[2370], lumberyards[2370]}), .right({trees[2372], lumberyards[2372]}), .bottom_left({trees[2420], lumberyards[2420]}), .bottom({trees[2421], lumberyards[2421]}), .bottom_right({trees[2422], lumberyards[2422]}), .init(2'b01), .state({trees[2371], lumberyards[2371]}));
acre acre_47_22 (.clk(clk), .en(en), .top_left({trees[2321], lumberyards[2321]}), .top({trees[2322], lumberyards[2322]}), .top_right({trees[2323], lumberyards[2323]}), .left({trees[2371], lumberyards[2371]}), .right({trees[2373], lumberyards[2373]}), .bottom_left({trees[2421], lumberyards[2421]}), .bottom({trees[2422], lumberyards[2422]}), .bottom_right({trees[2423], lumberyards[2423]}), .init(2'b10), .state({trees[2372], lumberyards[2372]}));
acre acre_47_23 (.clk(clk), .en(en), .top_left({trees[2322], lumberyards[2322]}), .top({trees[2323], lumberyards[2323]}), .top_right({trees[2324], lumberyards[2324]}), .left({trees[2372], lumberyards[2372]}), .right({trees[2374], lumberyards[2374]}), .bottom_left({trees[2422], lumberyards[2422]}), .bottom({trees[2423], lumberyards[2423]}), .bottom_right({trees[2424], lumberyards[2424]}), .init(2'b01), .state({trees[2373], lumberyards[2373]}));
acre acre_47_24 (.clk(clk), .en(en), .top_left({trees[2323], lumberyards[2323]}), .top({trees[2324], lumberyards[2324]}), .top_right({trees[2325], lumberyards[2325]}), .left({trees[2373], lumberyards[2373]}), .right({trees[2375], lumberyards[2375]}), .bottom_left({trees[2423], lumberyards[2423]}), .bottom({trees[2424], lumberyards[2424]}), .bottom_right({trees[2425], lumberyards[2425]}), .init(2'b00), .state({trees[2374], lumberyards[2374]}));
acre acre_47_25 (.clk(clk), .en(en), .top_left({trees[2324], lumberyards[2324]}), .top({trees[2325], lumberyards[2325]}), .top_right({trees[2326], lumberyards[2326]}), .left({trees[2374], lumberyards[2374]}), .right({trees[2376], lumberyards[2376]}), .bottom_left({trees[2424], lumberyards[2424]}), .bottom({trees[2425], lumberyards[2425]}), .bottom_right({trees[2426], lumberyards[2426]}), .init(2'b00), .state({trees[2375], lumberyards[2375]}));
acre acre_47_26 (.clk(clk), .en(en), .top_left({trees[2325], lumberyards[2325]}), .top({trees[2326], lumberyards[2326]}), .top_right({trees[2327], lumberyards[2327]}), .left({trees[2375], lumberyards[2375]}), .right({trees[2377], lumberyards[2377]}), .bottom_left({trees[2425], lumberyards[2425]}), .bottom({trees[2426], lumberyards[2426]}), .bottom_right({trees[2427], lumberyards[2427]}), .init(2'b10), .state({trees[2376], lumberyards[2376]}));
acre acre_47_27 (.clk(clk), .en(en), .top_left({trees[2326], lumberyards[2326]}), .top({trees[2327], lumberyards[2327]}), .top_right({trees[2328], lumberyards[2328]}), .left({trees[2376], lumberyards[2376]}), .right({trees[2378], lumberyards[2378]}), .bottom_left({trees[2426], lumberyards[2426]}), .bottom({trees[2427], lumberyards[2427]}), .bottom_right({trees[2428], lumberyards[2428]}), .init(2'b10), .state({trees[2377], lumberyards[2377]}));
acre acre_47_28 (.clk(clk), .en(en), .top_left({trees[2327], lumberyards[2327]}), .top({trees[2328], lumberyards[2328]}), .top_right({trees[2329], lumberyards[2329]}), .left({trees[2377], lumberyards[2377]}), .right({trees[2379], lumberyards[2379]}), .bottom_left({trees[2427], lumberyards[2427]}), .bottom({trees[2428], lumberyards[2428]}), .bottom_right({trees[2429], lumberyards[2429]}), .init(2'b00), .state({trees[2378], lumberyards[2378]}));
acre acre_47_29 (.clk(clk), .en(en), .top_left({trees[2328], lumberyards[2328]}), .top({trees[2329], lumberyards[2329]}), .top_right({trees[2330], lumberyards[2330]}), .left({trees[2378], lumberyards[2378]}), .right({trees[2380], lumberyards[2380]}), .bottom_left({trees[2428], lumberyards[2428]}), .bottom({trees[2429], lumberyards[2429]}), .bottom_right({trees[2430], lumberyards[2430]}), .init(2'b10), .state({trees[2379], lumberyards[2379]}));
acre acre_47_30 (.clk(clk), .en(en), .top_left({trees[2329], lumberyards[2329]}), .top({trees[2330], lumberyards[2330]}), .top_right({trees[2331], lumberyards[2331]}), .left({trees[2379], lumberyards[2379]}), .right({trees[2381], lumberyards[2381]}), .bottom_left({trees[2429], lumberyards[2429]}), .bottom({trees[2430], lumberyards[2430]}), .bottom_right({trees[2431], lumberyards[2431]}), .init(2'b10), .state({trees[2380], lumberyards[2380]}));
acre acre_47_31 (.clk(clk), .en(en), .top_left({trees[2330], lumberyards[2330]}), .top({trees[2331], lumberyards[2331]}), .top_right({trees[2332], lumberyards[2332]}), .left({trees[2380], lumberyards[2380]}), .right({trees[2382], lumberyards[2382]}), .bottom_left({trees[2430], lumberyards[2430]}), .bottom({trees[2431], lumberyards[2431]}), .bottom_right({trees[2432], lumberyards[2432]}), .init(2'b00), .state({trees[2381], lumberyards[2381]}));
acre acre_47_32 (.clk(clk), .en(en), .top_left({trees[2331], lumberyards[2331]}), .top({trees[2332], lumberyards[2332]}), .top_right({trees[2333], lumberyards[2333]}), .left({trees[2381], lumberyards[2381]}), .right({trees[2383], lumberyards[2383]}), .bottom_left({trees[2431], lumberyards[2431]}), .bottom({trees[2432], lumberyards[2432]}), .bottom_right({trees[2433], lumberyards[2433]}), .init(2'b00), .state({trees[2382], lumberyards[2382]}));
acre acre_47_33 (.clk(clk), .en(en), .top_left({trees[2332], lumberyards[2332]}), .top({trees[2333], lumberyards[2333]}), .top_right({trees[2334], lumberyards[2334]}), .left({trees[2382], lumberyards[2382]}), .right({trees[2384], lumberyards[2384]}), .bottom_left({trees[2432], lumberyards[2432]}), .bottom({trees[2433], lumberyards[2433]}), .bottom_right({trees[2434], lumberyards[2434]}), .init(2'b00), .state({trees[2383], lumberyards[2383]}));
acre acre_47_34 (.clk(clk), .en(en), .top_left({trees[2333], lumberyards[2333]}), .top({trees[2334], lumberyards[2334]}), .top_right({trees[2335], lumberyards[2335]}), .left({trees[2383], lumberyards[2383]}), .right({trees[2385], lumberyards[2385]}), .bottom_left({trees[2433], lumberyards[2433]}), .bottom({trees[2434], lumberyards[2434]}), .bottom_right({trees[2435], lumberyards[2435]}), .init(2'b00), .state({trees[2384], lumberyards[2384]}));
acre acre_47_35 (.clk(clk), .en(en), .top_left({trees[2334], lumberyards[2334]}), .top({trees[2335], lumberyards[2335]}), .top_right({trees[2336], lumberyards[2336]}), .left({trees[2384], lumberyards[2384]}), .right({trees[2386], lumberyards[2386]}), .bottom_left({trees[2434], lumberyards[2434]}), .bottom({trees[2435], lumberyards[2435]}), .bottom_right({trees[2436], lumberyards[2436]}), .init(2'b10), .state({trees[2385], lumberyards[2385]}));
acre acre_47_36 (.clk(clk), .en(en), .top_left({trees[2335], lumberyards[2335]}), .top({trees[2336], lumberyards[2336]}), .top_right({trees[2337], lumberyards[2337]}), .left({trees[2385], lumberyards[2385]}), .right({trees[2387], lumberyards[2387]}), .bottom_left({trees[2435], lumberyards[2435]}), .bottom({trees[2436], lumberyards[2436]}), .bottom_right({trees[2437], lumberyards[2437]}), .init(2'b00), .state({trees[2386], lumberyards[2386]}));
acre acre_47_37 (.clk(clk), .en(en), .top_left({trees[2336], lumberyards[2336]}), .top({trees[2337], lumberyards[2337]}), .top_right({trees[2338], lumberyards[2338]}), .left({trees[2386], lumberyards[2386]}), .right({trees[2388], lumberyards[2388]}), .bottom_left({trees[2436], lumberyards[2436]}), .bottom({trees[2437], lumberyards[2437]}), .bottom_right({trees[2438], lumberyards[2438]}), .init(2'b10), .state({trees[2387], lumberyards[2387]}));
acre acre_47_38 (.clk(clk), .en(en), .top_left({trees[2337], lumberyards[2337]}), .top({trees[2338], lumberyards[2338]}), .top_right({trees[2339], lumberyards[2339]}), .left({trees[2387], lumberyards[2387]}), .right({trees[2389], lumberyards[2389]}), .bottom_left({trees[2437], lumberyards[2437]}), .bottom({trees[2438], lumberyards[2438]}), .bottom_right({trees[2439], lumberyards[2439]}), .init(2'b00), .state({trees[2388], lumberyards[2388]}));
acre acre_47_39 (.clk(clk), .en(en), .top_left({trees[2338], lumberyards[2338]}), .top({trees[2339], lumberyards[2339]}), .top_right({trees[2340], lumberyards[2340]}), .left({trees[2388], lumberyards[2388]}), .right({trees[2390], lumberyards[2390]}), .bottom_left({trees[2438], lumberyards[2438]}), .bottom({trees[2439], lumberyards[2439]}), .bottom_right({trees[2440], lumberyards[2440]}), .init(2'b00), .state({trees[2389], lumberyards[2389]}));
acre acre_47_40 (.clk(clk), .en(en), .top_left({trees[2339], lumberyards[2339]}), .top({trees[2340], lumberyards[2340]}), .top_right({trees[2341], lumberyards[2341]}), .left({trees[2389], lumberyards[2389]}), .right({trees[2391], lumberyards[2391]}), .bottom_left({trees[2439], lumberyards[2439]}), .bottom({trees[2440], lumberyards[2440]}), .bottom_right({trees[2441], lumberyards[2441]}), .init(2'b00), .state({trees[2390], lumberyards[2390]}));
acre acre_47_41 (.clk(clk), .en(en), .top_left({trees[2340], lumberyards[2340]}), .top({trees[2341], lumberyards[2341]}), .top_right({trees[2342], lumberyards[2342]}), .left({trees[2390], lumberyards[2390]}), .right({trees[2392], lumberyards[2392]}), .bottom_left({trees[2440], lumberyards[2440]}), .bottom({trees[2441], lumberyards[2441]}), .bottom_right({trees[2442], lumberyards[2442]}), .init(2'b01), .state({trees[2391], lumberyards[2391]}));
acre acre_47_42 (.clk(clk), .en(en), .top_left({trees[2341], lumberyards[2341]}), .top({trees[2342], lumberyards[2342]}), .top_right({trees[2343], lumberyards[2343]}), .left({trees[2391], lumberyards[2391]}), .right({trees[2393], lumberyards[2393]}), .bottom_left({trees[2441], lumberyards[2441]}), .bottom({trees[2442], lumberyards[2442]}), .bottom_right({trees[2443], lumberyards[2443]}), .init(2'b00), .state({trees[2392], lumberyards[2392]}));
acre acre_47_43 (.clk(clk), .en(en), .top_left({trees[2342], lumberyards[2342]}), .top({trees[2343], lumberyards[2343]}), .top_right({trees[2344], lumberyards[2344]}), .left({trees[2392], lumberyards[2392]}), .right({trees[2394], lumberyards[2394]}), .bottom_left({trees[2442], lumberyards[2442]}), .bottom({trees[2443], lumberyards[2443]}), .bottom_right({trees[2444], lumberyards[2444]}), .init(2'b00), .state({trees[2393], lumberyards[2393]}));
acre acre_47_44 (.clk(clk), .en(en), .top_left({trees[2343], lumberyards[2343]}), .top({trees[2344], lumberyards[2344]}), .top_right({trees[2345], lumberyards[2345]}), .left({trees[2393], lumberyards[2393]}), .right({trees[2395], lumberyards[2395]}), .bottom_left({trees[2443], lumberyards[2443]}), .bottom({trees[2444], lumberyards[2444]}), .bottom_right({trees[2445], lumberyards[2445]}), .init(2'b01), .state({trees[2394], lumberyards[2394]}));
acre acre_47_45 (.clk(clk), .en(en), .top_left({trees[2344], lumberyards[2344]}), .top({trees[2345], lumberyards[2345]}), .top_right({trees[2346], lumberyards[2346]}), .left({trees[2394], lumberyards[2394]}), .right({trees[2396], lumberyards[2396]}), .bottom_left({trees[2444], lumberyards[2444]}), .bottom({trees[2445], lumberyards[2445]}), .bottom_right({trees[2446], lumberyards[2446]}), .init(2'b00), .state({trees[2395], lumberyards[2395]}));
acre acre_47_46 (.clk(clk), .en(en), .top_left({trees[2345], lumberyards[2345]}), .top({trees[2346], lumberyards[2346]}), .top_right({trees[2347], lumberyards[2347]}), .left({trees[2395], lumberyards[2395]}), .right({trees[2397], lumberyards[2397]}), .bottom_left({trees[2445], lumberyards[2445]}), .bottom({trees[2446], lumberyards[2446]}), .bottom_right({trees[2447], lumberyards[2447]}), .init(2'b10), .state({trees[2396], lumberyards[2396]}));
acre acre_47_47 (.clk(clk), .en(en), .top_left({trees[2346], lumberyards[2346]}), .top({trees[2347], lumberyards[2347]}), .top_right({trees[2348], lumberyards[2348]}), .left({trees[2396], lumberyards[2396]}), .right({trees[2398], lumberyards[2398]}), .bottom_left({trees[2446], lumberyards[2446]}), .bottom({trees[2447], lumberyards[2447]}), .bottom_right({trees[2448], lumberyards[2448]}), .init(2'b10), .state({trees[2397], lumberyards[2397]}));
acre acre_47_48 (.clk(clk), .en(en), .top_left({trees[2347], lumberyards[2347]}), .top({trees[2348], lumberyards[2348]}), .top_right({trees[2349], lumberyards[2349]}), .left({trees[2397], lumberyards[2397]}), .right({trees[2399], lumberyards[2399]}), .bottom_left({trees[2447], lumberyards[2447]}), .bottom({trees[2448], lumberyards[2448]}), .bottom_right({trees[2449], lumberyards[2449]}), .init(2'b00), .state({trees[2398], lumberyards[2398]}));
acre acre_47_49 (.clk(clk), .en(en), .top_left({trees[2348], lumberyards[2348]}), .top({trees[2349], lumberyards[2349]}), .top_right(2'b0), .left({trees[2398], lumberyards[2398]}), .right(2'b0), .bottom_left({trees[2448], lumberyards[2448]}), .bottom({trees[2449], lumberyards[2449]}), .bottom_right(2'b0), .init(2'b00), .state({trees[2399], lumberyards[2399]}));
acre acre_48_0 (.clk(clk), .en(en), .top_left(2'b0), .top({trees[2350], lumberyards[2350]}), .top_right({trees[2351], lumberyards[2351]}), .left(2'b0), .right({trees[2401], lumberyards[2401]}), .bottom_left(2'b0), .bottom({trees[2450], lumberyards[2450]}), .bottom_right({trees[2451], lumberyards[2451]}), .init(2'b10), .state({trees[2400], lumberyards[2400]}));
acre acre_48_1 (.clk(clk), .en(en), .top_left({trees[2350], lumberyards[2350]}), .top({trees[2351], lumberyards[2351]}), .top_right({trees[2352], lumberyards[2352]}), .left({trees[2400], lumberyards[2400]}), .right({trees[2402], lumberyards[2402]}), .bottom_left({trees[2450], lumberyards[2450]}), .bottom({trees[2451], lumberyards[2451]}), .bottom_right({trees[2452], lumberyards[2452]}), .init(2'b00), .state({trees[2401], lumberyards[2401]}));
acre acre_48_2 (.clk(clk), .en(en), .top_left({trees[2351], lumberyards[2351]}), .top({trees[2352], lumberyards[2352]}), .top_right({trees[2353], lumberyards[2353]}), .left({trees[2401], lumberyards[2401]}), .right({trees[2403], lumberyards[2403]}), .bottom_left({trees[2451], lumberyards[2451]}), .bottom({trees[2452], lumberyards[2452]}), .bottom_right({trees[2453], lumberyards[2453]}), .init(2'b01), .state({trees[2402], lumberyards[2402]}));
acre acre_48_3 (.clk(clk), .en(en), .top_left({trees[2352], lumberyards[2352]}), .top({trees[2353], lumberyards[2353]}), .top_right({trees[2354], lumberyards[2354]}), .left({trees[2402], lumberyards[2402]}), .right({trees[2404], lumberyards[2404]}), .bottom_left({trees[2452], lumberyards[2452]}), .bottom({trees[2453], lumberyards[2453]}), .bottom_right({trees[2454], lumberyards[2454]}), .init(2'b01), .state({trees[2403], lumberyards[2403]}));
acre acre_48_4 (.clk(clk), .en(en), .top_left({trees[2353], lumberyards[2353]}), .top({trees[2354], lumberyards[2354]}), .top_right({trees[2355], lumberyards[2355]}), .left({trees[2403], lumberyards[2403]}), .right({trees[2405], lumberyards[2405]}), .bottom_left({trees[2453], lumberyards[2453]}), .bottom({trees[2454], lumberyards[2454]}), .bottom_right({trees[2455], lumberyards[2455]}), .init(2'b00), .state({trees[2404], lumberyards[2404]}));
acre acre_48_5 (.clk(clk), .en(en), .top_left({trees[2354], lumberyards[2354]}), .top({trees[2355], lumberyards[2355]}), .top_right({trees[2356], lumberyards[2356]}), .left({trees[2404], lumberyards[2404]}), .right({trees[2406], lumberyards[2406]}), .bottom_left({trees[2454], lumberyards[2454]}), .bottom({trees[2455], lumberyards[2455]}), .bottom_right({trees[2456], lumberyards[2456]}), .init(2'b00), .state({trees[2405], lumberyards[2405]}));
acre acre_48_6 (.clk(clk), .en(en), .top_left({trees[2355], lumberyards[2355]}), .top({trees[2356], lumberyards[2356]}), .top_right({trees[2357], lumberyards[2357]}), .left({trees[2405], lumberyards[2405]}), .right({trees[2407], lumberyards[2407]}), .bottom_left({trees[2455], lumberyards[2455]}), .bottom({trees[2456], lumberyards[2456]}), .bottom_right({trees[2457], lumberyards[2457]}), .init(2'b01), .state({trees[2406], lumberyards[2406]}));
acre acre_48_7 (.clk(clk), .en(en), .top_left({trees[2356], lumberyards[2356]}), .top({trees[2357], lumberyards[2357]}), .top_right({trees[2358], lumberyards[2358]}), .left({trees[2406], lumberyards[2406]}), .right({trees[2408], lumberyards[2408]}), .bottom_left({trees[2456], lumberyards[2456]}), .bottom({trees[2457], lumberyards[2457]}), .bottom_right({trees[2458], lumberyards[2458]}), .init(2'b00), .state({trees[2407], lumberyards[2407]}));
acre acre_48_8 (.clk(clk), .en(en), .top_left({trees[2357], lumberyards[2357]}), .top({trees[2358], lumberyards[2358]}), .top_right({trees[2359], lumberyards[2359]}), .left({trees[2407], lumberyards[2407]}), .right({trees[2409], lumberyards[2409]}), .bottom_left({trees[2457], lumberyards[2457]}), .bottom({trees[2458], lumberyards[2458]}), .bottom_right({trees[2459], lumberyards[2459]}), .init(2'b00), .state({trees[2408], lumberyards[2408]}));
acre acre_48_9 (.clk(clk), .en(en), .top_left({trees[2358], lumberyards[2358]}), .top({trees[2359], lumberyards[2359]}), .top_right({trees[2360], lumberyards[2360]}), .left({trees[2408], lumberyards[2408]}), .right({trees[2410], lumberyards[2410]}), .bottom_left({trees[2458], lumberyards[2458]}), .bottom({trees[2459], lumberyards[2459]}), .bottom_right({trees[2460], lumberyards[2460]}), .init(2'b10), .state({trees[2409], lumberyards[2409]}));
acre acre_48_10 (.clk(clk), .en(en), .top_left({trees[2359], lumberyards[2359]}), .top({trees[2360], lumberyards[2360]}), .top_right({trees[2361], lumberyards[2361]}), .left({trees[2409], lumberyards[2409]}), .right({trees[2411], lumberyards[2411]}), .bottom_left({trees[2459], lumberyards[2459]}), .bottom({trees[2460], lumberyards[2460]}), .bottom_right({trees[2461], lumberyards[2461]}), .init(2'b00), .state({trees[2410], lumberyards[2410]}));
acre acre_48_11 (.clk(clk), .en(en), .top_left({trees[2360], lumberyards[2360]}), .top({trees[2361], lumberyards[2361]}), .top_right({trees[2362], lumberyards[2362]}), .left({trees[2410], lumberyards[2410]}), .right({trees[2412], lumberyards[2412]}), .bottom_left({trees[2460], lumberyards[2460]}), .bottom({trees[2461], lumberyards[2461]}), .bottom_right({trees[2462], lumberyards[2462]}), .init(2'b00), .state({trees[2411], lumberyards[2411]}));
acre acre_48_12 (.clk(clk), .en(en), .top_left({trees[2361], lumberyards[2361]}), .top({trees[2362], lumberyards[2362]}), .top_right({trees[2363], lumberyards[2363]}), .left({trees[2411], lumberyards[2411]}), .right({trees[2413], lumberyards[2413]}), .bottom_left({trees[2461], lumberyards[2461]}), .bottom({trees[2462], lumberyards[2462]}), .bottom_right({trees[2463], lumberyards[2463]}), .init(2'b00), .state({trees[2412], lumberyards[2412]}));
acre acre_48_13 (.clk(clk), .en(en), .top_left({trees[2362], lumberyards[2362]}), .top({trees[2363], lumberyards[2363]}), .top_right({trees[2364], lumberyards[2364]}), .left({trees[2412], lumberyards[2412]}), .right({trees[2414], lumberyards[2414]}), .bottom_left({trees[2462], lumberyards[2462]}), .bottom({trees[2463], lumberyards[2463]}), .bottom_right({trees[2464], lumberyards[2464]}), .init(2'b10), .state({trees[2413], lumberyards[2413]}));
acre acre_48_14 (.clk(clk), .en(en), .top_left({trees[2363], lumberyards[2363]}), .top({trees[2364], lumberyards[2364]}), .top_right({trees[2365], lumberyards[2365]}), .left({trees[2413], lumberyards[2413]}), .right({trees[2415], lumberyards[2415]}), .bottom_left({trees[2463], lumberyards[2463]}), .bottom({trees[2464], lumberyards[2464]}), .bottom_right({trees[2465], lumberyards[2465]}), .init(2'b10), .state({trees[2414], lumberyards[2414]}));
acre acre_48_15 (.clk(clk), .en(en), .top_left({trees[2364], lumberyards[2364]}), .top({trees[2365], lumberyards[2365]}), .top_right({trees[2366], lumberyards[2366]}), .left({trees[2414], lumberyards[2414]}), .right({trees[2416], lumberyards[2416]}), .bottom_left({trees[2464], lumberyards[2464]}), .bottom({trees[2465], lumberyards[2465]}), .bottom_right({trees[2466], lumberyards[2466]}), .init(2'b00), .state({trees[2415], lumberyards[2415]}));
acre acre_48_16 (.clk(clk), .en(en), .top_left({trees[2365], lumberyards[2365]}), .top({trees[2366], lumberyards[2366]}), .top_right({trees[2367], lumberyards[2367]}), .left({trees[2415], lumberyards[2415]}), .right({trees[2417], lumberyards[2417]}), .bottom_left({trees[2465], lumberyards[2465]}), .bottom({trees[2466], lumberyards[2466]}), .bottom_right({trees[2467], lumberyards[2467]}), .init(2'b10), .state({trees[2416], lumberyards[2416]}));
acre acre_48_17 (.clk(clk), .en(en), .top_left({trees[2366], lumberyards[2366]}), .top({trees[2367], lumberyards[2367]}), .top_right({trees[2368], lumberyards[2368]}), .left({trees[2416], lumberyards[2416]}), .right({trees[2418], lumberyards[2418]}), .bottom_left({trees[2466], lumberyards[2466]}), .bottom({trees[2467], lumberyards[2467]}), .bottom_right({trees[2468], lumberyards[2468]}), .init(2'b00), .state({trees[2417], lumberyards[2417]}));
acre acre_48_18 (.clk(clk), .en(en), .top_left({trees[2367], lumberyards[2367]}), .top({trees[2368], lumberyards[2368]}), .top_right({trees[2369], lumberyards[2369]}), .left({trees[2417], lumberyards[2417]}), .right({trees[2419], lumberyards[2419]}), .bottom_left({trees[2467], lumberyards[2467]}), .bottom({trees[2468], lumberyards[2468]}), .bottom_right({trees[2469], lumberyards[2469]}), .init(2'b00), .state({trees[2418], lumberyards[2418]}));
acre acre_48_19 (.clk(clk), .en(en), .top_left({trees[2368], lumberyards[2368]}), .top({trees[2369], lumberyards[2369]}), .top_right({trees[2370], lumberyards[2370]}), .left({trees[2418], lumberyards[2418]}), .right({trees[2420], lumberyards[2420]}), .bottom_left({trees[2468], lumberyards[2468]}), .bottom({trees[2469], lumberyards[2469]}), .bottom_right({trees[2470], lumberyards[2470]}), .init(2'b01), .state({trees[2419], lumberyards[2419]}));
acre acre_48_20 (.clk(clk), .en(en), .top_left({trees[2369], lumberyards[2369]}), .top({trees[2370], lumberyards[2370]}), .top_right({trees[2371], lumberyards[2371]}), .left({trees[2419], lumberyards[2419]}), .right({trees[2421], lumberyards[2421]}), .bottom_left({trees[2469], lumberyards[2469]}), .bottom({trees[2470], lumberyards[2470]}), .bottom_right({trees[2471], lumberyards[2471]}), .init(2'b00), .state({trees[2420], lumberyards[2420]}));
acre acre_48_21 (.clk(clk), .en(en), .top_left({trees[2370], lumberyards[2370]}), .top({trees[2371], lumberyards[2371]}), .top_right({trees[2372], lumberyards[2372]}), .left({trees[2420], lumberyards[2420]}), .right({trees[2422], lumberyards[2422]}), .bottom_left({trees[2470], lumberyards[2470]}), .bottom({trees[2471], lumberyards[2471]}), .bottom_right({trees[2472], lumberyards[2472]}), .init(2'b00), .state({trees[2421], lumberyards[2421]}));
acre acre_48_22 (.clk(clk), .en(en), .top_left({trees[2371], lumberyards[2371]}), .top({trees[2372], lumberyards[2372]}), .top_right({trees[2373], lumberyards[2373]}), .left({trees[2421], lumberyards[2421]}), .right({trees[2423], lumberyards[2423]}), .bottom_left({trees[2471], lumberyards[2471]}), .bottom({trees[2472], lumberyards[2472]}), .bottom_right({trees[2473], lumberyards[2473]}), .init(2'b00), .state({trees[2422], lumberyards[2422]}));
acre acre_48_23 (.clk(clk), .en(en), .top_left({trees[2372], lumberyards[2372]}), .top({trees[2373], lumberyards[2373]}), .top_right({trees[2374], lumberyards[2374]}), .left({trees[2422], lumberyards[2422]}), .right({trees[2424], lumberyards[2424]}), .bottom_left({trees[2472], lumberyards[2472]}), .bottom({trees[2473], lumberyards[2473]}), .bottom_right({trees[2474], lumberyards[2474]}), .init(2'b00), .state({trees[2423], lumberyards[2423]}));
acre acre_48_24 (.clk(clk), .en(en), .top_left({trees[2373], lumberyards[2373]}), .top({trees[2374], lumberyards[2374]}), .top_right({trees[2375], lumberyards[2375]}), .left({trees[2423], lumberyards[2423]}), .right({trees[2425], lumberyards[2425]}), .bottom_left({trees[2473], lumberyards[2473]}), .bottom({trees[2474], lumberyards[2474]}), .bottom_right({trees[2475], lumberyards[2475]}), .init(2'b10), .state({trees[2424], lumberyards[2424]}));
acre acre_48_25 (.clk(clk), .en(en), .top_left({trees[2374], lumberyards[2374]}), .top({trees[2375], lumberyards[2375]}), .top_right({trees[2376], lumberyards[2376]}), .left({trees[2424], lumberyards[2424]}), .right({trees[2426], lumberyards[2426]}), .bottom_left({trees[2474], lumberyards[2474]}), .bottom({trees[2475], lumberyards[2475]}), .bottom_right({trees[2476], lumberyards[2476]}), .init(2'b00), .state({trees[2425], lumberyards[2425]}));
acre acre_48_26 (.clk(clk), .en(en), .top_left({trees[2375], lumberyards[2375]}), .top({trees[2376], lumberyards[2376]}), .top_right({trees[2377], lumberyards[2377]}), .left({trees[2425], lumberyards[2425]}), .right({trees[2427], lumberyards[2427]}), .bottom_left({trees[2475], lumberyards[2475]}), .bottom({trees[2476], lumberyards[2476]}), .bottom_right({trees[2477], lumberyards[2477]}), .init(2'b10), .state({trees[2426], lumberyards[2426]}));
acre acre_48_27 (.clk(clk), .en(en), .top_left({trees[2376], lumberyards[2376]}), .top({trees[2377], lumberyards[2377]}), .top_right({trees[2378], lumberyards[2378]}), .left({trees[2426], lumberyards[2426]}), .right({trees[2428], lumberyards[2428]}), .bottom_left({trees[2476], lumberyards[2476]}), .bottom({trees[2477], lumberyards[2477]}), .bottom_right({trees[2478], lumberyards[2478]}), .init(2'b00), .state({trees[2427], lumberyards[2427]}));
acre acre_48_28 (.clk(clk), .en(en), .top_left({trees[2377], lumberyards[2377]}), .top({trees[2378], lumberyards[2378]}), .top_right({trees[2379], lumberyards[2379]}), .left({trees[2427], lumberyards[2427]}), .right({trees[2429], lumberyards[2429]}), .bottom_left({trees[2477], lumberyards[2477]}), .bottom({trees[2478], lumberyards[2478]}), .bottom_right({trees[2479], lumberyards[2479]}), .init(2'b01), .state({trees[2428], lumberyards[2428]}));
acre acre_48_29 (.clk(clk), .en(en), .top_left({trees[2378], lumberyards[2378]}), .top({trees[2379], lumberyards[2379]}), .top_right({trees[2380], lumberyards[2380]}), .left({trees[2428], lumberyards[2428]}), .right({trees[2430], lumberyards[2430]}), .bottom_left({trees[2478], lumberyards[2478]}), .bottom({trees[2479], lumberyards[2479]}), .bottom_right({trees[2480], lumberyards[2480]}), .init(2'b10), .state({trees[2429], lumberyards[2429]}));
acre acre_48_30 (.clk(clk), .en(en), .top_left({trees[2379], lumberyards[2379]}), .top({trees[2380], lumberyards[2380]}), .top_right({trees[2381], lumberyards[2381]}), .left({trees[2429], lumberyards[2429]}), .right({trees[2431], lumberyards[2431]}), .bottom_left({trees[2479], lumberyards[2479]}), .bottom({trees[2480], lumberyards[2480]}), .bottom_right({trees[2481], lumberyards[2481]}), .init(2'b00), .state({trees[2430], lumberyards[2430]}));
acre acre_48_31 (.clk(clk), .en(en), .top_left({trees[2380], lumberyards[2380]}), .top({trees[2381], lumberyards[2381]}), .top_right({trees[2382], lumberyards[2382]}), .left({trees[2430], lumberyards[2430]}), .right({trees[2432], lumberyards[2432]}), .bottom_left({trees[2480], lumberyards[2480]}), .bottom({trees[2481], lumberyards[2481]}), .bottom_right({trees[2482], lumberyards[2482]}), .init(2'b00), .state({trees[2431], lumberyards[2431]}));
acre acre_48_32 (.clk(clk), .en(en), .top_left({trees[2381], lumberyards[2381]}), .top({trees[2382], lumberyards[2382]}), .top_right({trees[2383], lumberyards[2383]}), .left({trees[2431], lumberyards[2431]}), .right({trees[2433], lumberyards[2433]}), .bottom_left({trees[2481], lumberyards[2481]}), .bottom({trees[2482], lumberyards[2482]}), .bottom_right({trees[2483], lumberyards[2483]}), .init(2'b01), .state({trees[2432], lumberyards[2432]}));
acre acre_48_33 (.clk(clk), .en(en), .top_left({trees[2382], lumberyards[2382]}), .top({trees[2383], lumberyards[2383]}), .top_right({trees[2384], lumberyards[2384]}), .left({trees[2432], lumberyards[2432]}), .right({trees[2434], lumberyards[2434]}), .bottom_left({trees[2482], lumberyards[2482]}), .bottom({trees[2483], lumberyards[2483]}), .bottom_right({trees[2484], lumberyards[2484]}), .init(2'b00), .state({trees[2433], lumberyards[2433]}));
acre acre_48_34 (.clk(clk), .en(en), .top_left({trees[2383], lumberyards[2383]}), .top({trees[2384], lumberyards[2384]}), .top_right({trees[2385], lumberyards[2385]}), .left({trees[2433], lumberyards[2433]}), .right({trees[2435], lumberyards[2435]}), .bottom_left({trees[2483], lumberyards[2483]}), .bottom({trees[2484], lumberyards[2484]}), .bottom_right({trees[2485], lumberyards[2485]}), .init(2'b10), .state({trees[2434], lumberyards[2434]}));
acre acre_48_35 (.clk(clk), .en(en), .top_left({trees[2384], lumberyards[2384]}), .top({trees[2385], lumberyards[2385]}), .top_right({trees[2386], lumberyards[2386]}), .left({trees[2434], lumberyards[2434]}), .right({trees[2436], lumberyards[2436]}), .bottom_left({trees[2484], lumberyards[2484]}), .bottom({trees[2485], lumberyards[2485]}), .bottom_right({trees[2486], lumberyards[2486]}), .init(2'b10), .state({trees[2435], lumberyards[2435]}));
acre acre_48_36 (.clk(clk), .en(en), .top_left({trees[2385], lumberyards[2385]}), .top({trees[2386], lumberyards[2386]}), .top_right({trees[2387], lumberyards[2387]}), .left({trees[2435], lumberyards[2435]}), .right({trees[2437], lumberyards[2437]}), .bottom_left({trees[2485], lumberyards[2485]}), .bottom({trees[2486], lumberyards[2486]}), .bottom_right({trees[2487], lumberyards[2487]}), .init(2'b00), .state({trees[2436], lumberyards[2436]}));
acre acre_48_37 (.clk(clk), .en(en), .top_left({trees[2386], lumberyards[2386]}), .top({trees[2387], lumberyards[2387]}), .top_right({trees[2388], lumberyards[2388]}), .left({trees[2436], lumberyards[2436]}), .right({trees[2438], lumberyards[2438]}), .bottom_left({trees[2486], lumberyards[2486]}), .bottom({trees[2487], lumberyards[2487]}), .bottom_right({trees[2488], lumberyards[2488]}), .init(2'b00), .state({trees[2437], lumberyards[2437]}));
acre acre_48_38 (.clk(clk), .en(en), .top_left({trees[2387], lumberyards[2387]}), .top({trees[2388], lumberyards[2388]}), .top_right({trees[2389], lumberyards[2389]}), .left({trees[2437], lumberyards[2437]}), .right({trees[2439], lumberyards[2439]}), .bottom_left({trees[2487], lumberyards[2487]}), .bottom({trees[2488], lumberyards[2488]}), .bottom_right({trees[2489], lumberyards[2489]}), .init(2'b01), .state({trees[2438], lumberyards[2438]}));
acre acre_48_39 (.clk(clk), .en(en), .top_left({trees[2388], lumberyards[2388]}), .top({trees[2389], lumberyards[2389]}), .top_right({trees[2390], lumberyards[2390]}), .left({trees[2438], lumberyards[2438]}), .right({trees[2440], lumberyards[2440]}), .bottom_left({trees[2488], lumberyards[2488]}), .bottom({trees[2489], lumberyards[2489]}), .bottom_right({trees[2490], lumberyards[2490]}), .init(2'b00), .state({trees[2439], lumberyards[2439]}));
acre acre_48_40 (.clk(clk), .en(en), .top_left({trees[2389], lumberyards[2389]}), .top({trees[2390], lumberyards[2390]}), .top_right({trees[2391], lumberyards[2391]}), .left({trees[2439], lumberyards[2439]}), .right({trees[2441], lumberyards[2441]}), .bottom_left({trees[2489], lumberyards[2489]}), .bottom({trees[2490], lumberyards[2490]}), .bottom_right({trees[2491], lumberyards[2491]}), .init(2'b00), .state({trees[2440], lumberyards[2440]}));
acre acre_48_41 (.clk(clk), .en(en), .top_left({trees[2390], lumberyards[2390]}), .top({trees[2391], lumberyards[2391]}), .top_right({trees[2392], lumberyards[2392]}), .left({trees[2440], lumberyards[2440]}), .right({trees[2442], lumberyards[2442]}), .bottom_left({trees[2490], lumberyards[2490]}), .bottom({trees[2491], lumberyards[2491]}), .bottom_right({trees[2492], lumberyards[2492]}), .init(2'b01), .state({trees[2441], lumberyards[2441]}));
acre acre_48_42 (.clk(clk), .en(en), .top_left({trees[2391], lumberyards[2391]}), .top({trees[2392], lumberyards[2392]}), .top_right({trees[2393], lumberyards[2393]}), .left({trees[2441], lumberyards[2441]}), .right({trees[2443], lumberyards[2443]}), .bottom_left({trees[2491], lumberyards[2491]}), .bottom({trees[2492], lumberyards[2492]}), .bottom_right({trees[2493], lumberyards[2493]}), .init(2'b01), .state({trees[2442], lumberyards[2442]}));
acre acre_48_43 (.clk(clk), .en(en), .top_left({trees[2392], lumberyards[2392]}), .top({trees[2393], lumberyards[2393]}), .top_right({trees[2394], lumberyards[2394]}), .left({trees[2442], lumberyards[2442]}), .right({trees[2444], lumberyards[2444]}), .bottom_left({trees[2492], lumberyards[2492]}), .bottom({trees[2493], lumberyards[2493]}), .bottom_right({trees[2494], lumberyards[2494]}), .init(2'b01), .state({trees[2443], lumberyards[2443]}));
acre acre_48_44 (.clk(clk), .en(en), .top_left({trees[2393], lumberyards[2393]}), .top({trees[2394], lumberyards[2394]}), .top_right({trees[2395], lumberyards[2395]}), .left({trees[2443], lumberyards[2443]}), .right({trees[2445], lumberyards[2445]}), .bottom_left({trees[2493], lumberyards[2493]}), .bottom({trees[2494], lumberyards[2494]}), .bottom_right({trees[2495], lumberyards[2495]}), .init(2'b01), .state({trees[2444], lumberyards[2444]}));
acre acre_48_45 (.clk(clk), .en(en), .top_left({trees[2394], lumberyards[2394]}), .top({trees[2395], lumberyards[2395]}), .top_right({trees[2396], lumberyards[2396]}), .left({trees[2444], lumberyards[2444]}), .right({trees[2446], lumberyards[2446]}), .bottom_left({trees[2494], lumberyards[2494]}), .bottom({trees[2495], lumberyards[2495]}), .bottom_right({trees[2496], lumberyards[2496]}), .init(2'b00), .state({trees[2445], lumberyards[2445]}));
acre acre_48_46 (.clk(clk), .en(en), .top_left({trees[2395], lumberyards[2395]}), .top({trees[2396], lumberyards[2396]}), .top_right({trees[2397], lumberyards[2397]}), .left({trees[2445], lumberyards[2445]}), .right({trees[2447], lumberyards[2447]}), .bottom_left({trees[2495], lumberyards[2495]}), .bottom({trees[2496], lumberyards[2496]}), .bottom_right({trees[2497], lumberyards[2497]}), .init(2'b01), .state({trees[2446], lumberyards[2446]}));
acre acre_48_47 (.clk(clk), .en(en), .top_left({trees[2396], lumberyards[2396]}), .top({trees[2397], lumberyards[2397]}), .top_right({trees[2398], lumberyards[2398]}), .left({trees[2446], lumberyards[2446]}), .right({trees[2448], lumberyards[2448]}), .bottom_left({trees[2496], lumberyards[2496]}), .bottom({trees[2497], lumberyards[2497]}), .bottom_right({trees[2498], lumberyards[2498]}), .init(2'b00), .state({trees[2447], lumberyards[2447]}));
acre acre_48_48 (.clk(clk), .en(en), .top_left({trees[2397], lumberyards[2397]}), .top({trees[2398], lumberyards[2398]}), .top_right({trees[2399], lumberyards[2399]}), .left({trees[2447], lumberyards[2447]}), .right({trees[2449], lumberyards[2449]}), .bottom_left({trees[2497], lumberyards[2497]}), .bottom({trees[2498], lumberyards[2498]}), .bottom_right({trees[2499], lumberyards[2499]}), .init(2'b00), .state({trees[2448], lumberyards[2448]}));
acre acre_48_49 (.clk(clk), .en(en), .top_left({trees[2398], lumberyards[2398]}), .top({trees[2399], lumberyards[2399]}), .top_right(2'b0), .left({trees[2448], lumberyards[2448]}), .right(2'b0), .bottom_left({trees[2498], lumberyards[2498]}), .bottom({trees[2499], lumberyards[2499]}), .bottom_right(2'b0), .init(2'b00), .state({trees[2449], lumberyards[2449]}));
acre acre_49_0 (.clk(clk), .en(en), .top_left(2'b0), .top({trees[2400], lumberyards[2400]}), .top_right({trees[2401], lumberyards[2401]}), .left(2'b0), .right({trees[2451], lumberyards[2451]}), .bottom_left(2'b0), .bottom(2'b0), .bottom_right(2'b0), .init(2'b00), .state({trees[2450], lumberyards[2450]}));
acre acre_49_1 (.clk(clk), .en(en), .top_left({trees[2400], lumberyards[2400]}), .top({trees[2401], lumberyards[2401]}), .top_right({trees[2402], lumberyards[2402]}), .left({trees[2450], lumberyards[2450]}), .right({trees[2452], lumberyards[2452]}), .bottom_left(2'b0), .bottom(2'b0), .bottom_right(2'b0), .init(2'b10), .state({trees[2451], lumberyards[2451]}));
acre acre_49_2 (.clk(clk), .en(en), .top_left({trees[2401], lumberyards[2401]}), .top({trees[2402], lumberyards[2402]}), .top_right({trees[2403], lumberyards[2403]}), .left({trees[2451], lumberyards[2451]}), .right({trees[2453], lumberyards[2453]}), .bottom_left(2'b0), .bottom(2'b0), .bottom_right(2'b0), .init(2'b10), .state({trees[2452], lumberyards[2452]}));
acre acre_49_3 (.clk(clk), .en(en), .top_left({trees[2402], lumberyards[2402]}), .top({trees[2403], lumberyards[2403]}), .top_right({trees[2404], lumberyards[2404]}), .left({trees[2452], lumberyards[2452]}), .right({trees[2454], lumberyards[2454]}), .bottom_left(2'b0), .bottom(2'b0), .bottom_right(2'b0), .init(2'b00), .state({trees[2453], lumberyards[2453]}));
acre acre_49_4 (.clk(clk), .en(en), .top_left({trees[2403], lumberyards[2403]}), .top({trees[2404], lumberyards[2404]}), .top_right({trees[2405], lumberyards[2405]}), .left({trees[2453], lumberyards[2453]}), .right({trees[2455], lumberyards[2455]}), .bottom_left(2'b0), .bottom(2'b0), .bottom_right(2'b0), .init(2'b00), .state({trees[2454], lumberyards[2454]}));
acre acre_49_5 (.clk(clk), .en(en), .top_left({trees[2404], lumberyards[2404]}), .top({trees[2405], lumberyards[2405]}), .top_right({trees[2406], lumberyards[2406]}), .left({trees[2454], lumberyards[2454]}), .right({trees[2456], lumberyards[2456]}), .bottom_left(2'b0), .bottom(2'b0), .bottom_right(2'b0), .init(2'b10), .state({trees[2455], lumberyards[2455]}));
acre acre_49_6 (.clk(clk), .en(en), .top_left({trees[2405], lumberyards[2405]}), .top({trees[2406], lumberyards[2406]}), .top_right({trees[2407], lumberyards[2407]}), .left({trees[2455], lumberyards[2455]}), .right({trees[2457], lumberyards[2457]}), .bottom_left(2'b0), .bottom(2'b0), .bottom_right(2'b0), .init(2'b00), .state({trees[2456], lumberyards[2456]}));
acre acre_49_7 (.clk(clk), .en(en), .top_left({trees[2406], lumberyards[2406]}), .top({trees[2407], lumberyards[2407]}), .top_right({trees[2408], lumberyards[2408]}), .left({trees[2456], lumberyards[2456]}), .right({trees[2458], lumberyards[2458]}), .bottom_left(2'b0), .bottom(2'b0), .bottom_right(2'b0), .init(2'b10), .state({trees[2457], lumberyards[2457]}));
acre acre_49_8 (.clk(clk), .en(en), .top_left({trees[2407], lumberyards[2407]}), .top({trees[2408], lumberyards[2408]}), .top_right({trees[2409], lumberyards[2409]}), .left({trees[2457], lumberyards[2457]}), .right({trees[2459], lumberyards[2459]}), .bottom_left(2'b0), .bottom(2'b0), .bottom_right(2'b0), .init(2'b00), .state({trees[2458], lumberyards[2458]}));
acre acre_49_9 (.clk(clk), .en(en), .top_left({trees[2408], lumberyards[2408]}), .top({trees[2409], lumberyards[2409]}), .top_right({trees[2410], lumberyards[2410]}), .left({trees[2458], lumberyards[2458]}), .right({trees[2460], lumberyards[2460]}), .bottom_left(2'b0), .bottom(2'b0), .bottom_right(2'b0), .init(2'b00), .state({trees[2459], lumberyards[2459]}));
acre acre_49_10 (.clk(clk), .en(en), .top_left({trees[2409], lumberyards[2409]}), .top({trees[2410], lumberyards[2410]}), .top_right({trees[2411], lumberyards[2411]}), .left({trees[2459], lumberyards[2459]}), .right({trees[2461], lumberyards[2461]}), .bottom_left(2'b0), .bottom(2'b0), .bottom_right(2'b0), .init(2'b00), .state({trees[2460], lumberyards[2460]}));
acre acre_49_11 (.clk(clk), .en(en), .top_left({trees[2410], lumberyards[2410]}), .top({trees[2411], lumberyards[2411]}), .top_right({trees[2412], lumberyards[2412]}), .left({trees[2460], lumberyards[2460]}), .right({trees[2462], lumberyards[2462]}), .bottom_left(2'b0), .bottom(2'b0), .bottom_right(2'b0), .init(2'b10), .state({trees[2461], lumberyards[2461]}));
acre acre_49_12 (.clk(clk), .en(en), .top_left({trees[2411], lumberyards[2411]}), .top({trees[2412], lumberyards[2412]}), .top_right({trees[2413], lumberyards[2413]}), .left({trees[2461], lumberyards[2461]}), .right({trees[2463], lumberyards[2463]}), .bottom_left(2'b0), .bottom(2'b0), .bottom_right(2'b0), .init(2'b01), .state({trees[2462], lumberyards[2462]}));
acre acre_49_13 (.clk(clk), .en(en), .top_left({trees[2412], lumberyards[2412]}), .top({trees[2413], lumberyards[2413]}), .top_right({trees[2414], lumberyards[2414]}), .left({trees[2462], lumberyards[2462]}), .right({trees[2464], lumberyards[2464]}), .bottom_left(2'b0), .bottom(2'b0), .bottom_right(2'b0), .init(2'b10), .state({trees[2463], lumberyards[2463]}));
acre acre_49_14 (.clk(clk), .en(en), .top_left({trees[2413], lumberyards[2413]}), .top({trees[2414], lumberyards[2414]}), .top_right({trees[2415], lumberyards[2415]}), .left({trees[2463], lumberyards[2463]}), .right({trees[2465], lumberyards[2465]}), .bottom_left(2'b0), .bottom(2'b0), .bottom_right(2'b0), .init(2'b01), .state({trees[2464], lumberyards[2464]}));
acre acre_49_15 (.clk(clk), .en(en), .top_left({trees[2414], lumberyards[2414]}), .top({trees[2415], lumberyards[2415]}), .top_right({trees[2416], lumberyards[2416]}), .left({trees[2464], lumberyards[2464]}), .right({trees[2466], lumberyards[2466]}), .bottom_left(2'b0), .bottom(2'b0), .bottom_right(2'b0), .init(2'b00), .state({trees[2465], lumberyards[2465]}));
acre acre_49_16 (.clk(clk), .en(en), .top_left({trees[2415], lumberyards[2415]}), .top({trees[2416], lumberyards[2416]}), .top_right({trees[2417], lumberyards[2417]}), .left({trees[2465], lumberyards[2465]}), .right({trees[2467], lumberyards[2467]}), .bottom_left(2'b0), .bottom(2'b0), .bottom_right(2'b0), .init(2'b10), .state({trees[2466], lumberyards[2466]}));
acre acre_49_17 (.clk(clk), .en(en), .top_left({trees[2416], lumberyards[2416]}), .top({trees[2417], lumberyards[2417]}), .top_right({trees[2418], lumberyards[2418]}), .left({trees[2466], lumberyards[2466]}), .right({trees[2468], lumberyards[2468]}), .bottom_left(2'b0), .bottom(2'b0), .bottom_right(2'b0), .init(2'b10), .state({trees[2467], lumberyards[2467]}));
acre acre_49_18 (.clk(clk), .en(en), .top_left({trees[2417], lumberyards[2417]}), .top({trees[2418], lumberyards[2418]}), .top_right({trees[2419], lumberyards[2419]}), .left({trees[2467], lumberyards[2467]}), .right({trees[2469], lumberyards[2469]}), .bottom_left(2'b0), .bottom(2'b0), .bottom_right(2'b0), .init(2'b10), .state({trees[2468], lumberyards[2468]}));
acre acre_49_19 (.clk(clk), .en(en), .top_left({trees[2418], lumberyards[2418]}), .top({trees[2419], lumberyards[2419]}), .top_right({trees[2420], lumberyards[2420]}), .left({trees[2468], lumberyards[2468]}), .right({trees[2470], lumberyards[2470]}), .bottom_left(2'b0), .bottom(2'b0), .bottom_right(2'b0), .init(2'b01), .state({trees[2469], lumberyards[2469]}));
acre acre_49_20 (.clk(clk), .en(en), .top_left({trees[2419], lumberyards[2419]}), .top({trees[2420], lumberyards[2420]}), .top_right({trees[2421], lumberyards[2421]}), .left({trees[2469], lumberyards[2469]}), .right({trees[2471], lumberyards[2471]}), .bottom_left(2'b0), .bottom(2'b0), .bottom_right(2'b0), .init(2'b00), .state({trees[2470], lumberyards[2470]}));
acre acre_49_21 (.clk(clk), .en(en), .top_left({trees[2420], lumberyards[2420]}), .top({trees[2421], lumberyards[2421]}), .top_right({trees[2422], lumberyards[2422]}), .left({trees[2470], lumberyards[2470]}), .right({trees[2472], lumberyards[2472]}), .bottom_left(2'b0), .bottom(2'b0), .bottom_right(2'b0), .init(2'b00), .state({trees[2471], lumberyards[2471]}));
acre acre_49_22 (.clk(clk), .en(en), .top_left({trees[2421], lumberyards[2421]}), .top({trees[2422], lumberyards[2422]}), .top_right({trees[2423], lumberyards[2423]}), .left({trees[2471], lumberyards[2471]}), .right({trees[2473], lumberyards[2473]}), .bottom_left(2'b0), .bottom(2'b0), .bottom_right(2'b0), .init(2'b00), .state({trees[2472], lumberyards[2472]}));
acre acre_49_23 (.clk(clk), .en(en), .top_left({trees[2422], lumberyards[2422]}), .top({trees[2423], lumberyards[2423]}), .top_right({trees[2424], lumberyards[2424]}), .left({trees[2472], lumberyards[2472]}), .right({trees[2474], lumberyards[2474]}), .bottom_left(2'b0), .bottom(2'b0), .bottom_right(2'b0), .init(2'b00), .state({trees[2473], lumberyards[2473]}));
acre acre_49_24 (.clk(clk), .en(en), .top_left({trees[2423], lumberyards[2423]}), .top({trees[2424], lumberyards[2424]}), .top_right({trees[2425], lumberyards[2425]}), .left({trees[2473], lumberyards[2473]}), .right({trees[2475], lumberyards[2475]}), .bottom_left(2'b0), .bottom(2'b0), .bottom_right(2'b0), .init(2'b00), .state({trees[2474], lumberyards[2474]}));
acre acre_49_25 (.clk(clk), .en(en), .top_left({trees[2424], lumberyards[2424]}), .top({trees[2425], lumberyards[2425]}), .top_right({trees[2426], lumberyards[2426]}), .left({trees[2474], lumberyards[2474]}), .right({trees[2476], lumberyards[2476]}), .bottom_left(2'b0), .bottom(2'b0), .bottom_right(2'b0), .init(2'b00), .state({trees[2475], lumberyards[2475]}));
acre acre_49_26 (.clk(clk), .en(en), .top_left({trees[2425], lumberyards[2425]}), .top({trees[2426], lumberyards[2426]}), .top_right({trees[2427], lumberyards[2427]}), .left({trees[2475], lumberyards[2475]}), .right({trees[2477], lumberyards[2477]}), .bottom_left(2'b0), .bottom(2'b0), .bottom_right(2'b0), .init(2'b10), .state({trees[2476], lumberyards[2476]}));
acre acre_49_27 (.clk(clk), .en(en), .top_left({trees[2426], lumberyards[2426]}), .top({trees[2427], lumberyards[2427]}), .top_right({trees[2428], lumberyards[2428]}), .left({trees[2476], lumberyards[2476]}), .right({trees[2478], lumberyards[2478]}), .bottom_left(2'b0), .bottom(2'b0), .bottom_right(2'b0), .init(2'b00), .state({trees[2477], lumberyards[2477]}));
acre acre_49_28 (.clk(clk), .en(en), .top_left({trees[2427], lumberyards[2427]}), .top({trees[2428], lumberyards[2428]}), .top_right({trees[2429], lumberyards[2429]}), .left({trees[2477], lumberyards[2477]}), .right({trees[2479], lumberyards[2479]}), .bottom_left(2'b0), .bottom(2'b0), .bottom_right(2'b0), .init(2'b00), .state({trees[2478], lumberyards[2478]}));
acre acre_49_29 (.clk(clk), .en(en), .top_left({trees[2428], lumberyards[2428]}), .top({trees[2429], lumberyards[2429]}), .top_right({trees[2430], lumberyards[2430]}), .left({trees[2478], lumberyards[2478]}), .right({trees[2480], lumberyards[2480]}), .bottom_left(2'b0), .bottom(2'b0), .bottom_right(2'b0), .init(2'b00), .state({trees[2479], lumberyards[2479]}));
acre acre_49_30 (.clk(clk), .en(en), .top_left({trees[2429], lumberyards[2429]}), .top({trees[2430], lumberyards[2430]}), .top_right({trees[2431], lumberyards[2431]}), .left({trees[2479], lumberyards[2479]}), .right({trees[2481], lumberyards[2481]}), .bottom_left(2'b0), .bottom(2'b0), .bottom_right(2'b0), .init(2'b00), .state({trees[2480], lumberyards[2480]}));
acre acre_49_31 (.clk(clk), .en(en), .top_left({trees[2430], lumberyards[2430]}), .top({trees[2431], lumberyards[2431]}), .top_right({trees[2432], lumberyards[2432]}), .left({trees[2480], lumberyards[2480]}), .right({trees[2482], lumberyards[2482]}), .bottom_left(2'b0), .bottom(2'b0), .bottom_right(2'b0), .init(2'b00), .state({trees[2481], lumberyards[2481]}));
acre acre_49_32 (.clk(clk), .en(en), .top_left({trees[2431], lumberyards[2431]}), .top({trees[2432], lumberyards[2432]}), .top_right({trees[2433], lumberyards[2433]}), .left({trees[2481], lumberyards[2481]}), .right({trees[2483], lumberyards[2483]}), .bottom_left(2'b0), .bottom(2'b0), .bottom_right(2'b0), .init(2'b00), .state({trees[2482], lumberyards[2482]}));
acre acre_49_33 (.clk(clk), .en(en), .top_left({trees[2432], lumberyards[2432]}), .top({trees[2433], lumberyards[2433]}), .top_right({trees[2434], lumberyards[2434]}), .left({trees[2482], lumberyards[2482]}), .right({trees[2484], lumberyards[2484]}), .bottom_left(2'b0), .bottom(2'b0), .bottom_right(2'b0), .init(2'b01), .state({trees[2483], lumberyards[2483]}));
acre acre_49_34 (.clk(clk), .en(en), .top_left({trees[2433], lumberyards[2433]}), .top({trees[2434], lumberyards[2434]}), .top_right({trees[2435], lumberyards[2435]}), .left({trees[2483], lumberyards[2483]}), .right({trees[2485], lumberyards[2485]}), .bottom_left(2'b0), .bottom(2'b0), .bottom_right(2'b0), .init(2'b00), .state({trees[2484], lumberyards[2484]}));
acre acre_49_35 (.clk(clk), .en(en), .top_left({trees[2434], lumberyards[2434]}), .top({trees[2435], lumberyards[2435]}), .top_right({trees[2436], lumberyards[2436]}), .left({trees[2484], lumberyards[2484]}), .right({trees[2486], lumberyards[2486]}), .bottom_left(2'b0), .bottom(2'b0), .bottom_right(2'b0), .init(2'b10), .state({trees[2485], lumberyards[2485]}));
acre acre_49_36 (.clk(clk), .en(en), .top_left({trees[2435], lumberyards[2435]}), .top({trees[2436], lumberyards[2436]}), .top_right({trees[2437], lumberyards[2437]}), .left({trees[2485], lumberyards[2485]}), .right({trees[2487], lumberyards[2487]}), .bottom_left(2'b0), .bottom(2'b0), .bottom_right(2'b0), .init(2'b00), .state({trees[2486], lumberyards[2486]}));
acre acre_49_37 (.clk(clk), .en(en), .top_left({trees[2436], lumberyards[2436]}), .top({trees[2437], lumberyards[2437]}), .top_right({trees[2438], lumberyards[2438]}), .left({trees[2486], lumberyards[2486]}), .right({trees[2488], lumberyards[2488]}), .bottom_left(2'b0), .bottom(2'b0), .bottom_right(2'b0), .init(2'b00), .state({trees[2487], lumberyards[2487]}));
acre acre_49_38 (.clk(clk), .en(en), .top_left({trees[2437], lumberyards[2437]}), .top({trees[2438], lumberyards[2438]}), .top_right({trees[2439], lumberyards[2439]}), .left({trees[2487], lumberyards[2487]}), .right({trees[2489], lumberyards[2489]}), .bottom_left(2'b0), .bottom(2'b0), .bottom_right(2'b0), .init(2'b00), .state({trees[2488], lumberyards[2488]}));
acre acre_49_39 (.clk(clk), .en(en), .top_left({trees[2438], lumberyards[2438]}), .top({trees[2439], lumberyards[2439]}), .top_right({trees[2440], lumberyards[2440]}), .left({trees[2488], lumberyards[2488]}), .right({trees[2490], lumberyards[2490]}), .bottom_left(2'b0), .bottom(2'b0), .bottom_right(2'b0), .init(2'b00), .state({trees[2489], lumberyards[2489]}));
acre acre_49_40 (.clk(clk), .en(en), .top_left({trees[2439], lumberyards[2439]}), .top({trees[2440], lumberyards[2440]}), .top_right({trees[2441], lumberyards[2441]}), .left({trees[2489], lumberyards[2489]}), .right({trees[2491], lumberyards[2491]}), .bottom_left(2'b0), .bottom(2'b0), .bottom_right(2'b0), .init(2'b00), .state({trees[2490], lumberyards[2490]}));
acre acre_49_41 (.clk(clk), .en(en), .top_left({trees[2440], lumberyards[2440]}), .top({trees[2441], lumberyards[2441]}), .top_right({trees[2442], lumberyards[2442]}), .left({trees[2490], lumberyards[2490]}), .right({trees[2492], lumberyards[2492]}), .bottom_left(2'b0), .bottom(2'b0), .bottom_right(2'b0), .init(2'b10), .state({trees[2491], lumberyards[2491]}));
acre acre_49_42 (.clk(clk), .en(en), .top_left({trees[2441], lumberyards[2441]}), .top({trees[2442], lumberyards[2442]}), .top_right({trees[2443], lumberyards[2443]}), .left({trees[2491], lumberyards[2491]}), .right({trees[2493], lumberyards[2493]}), .bottom_left(2'b0), .bottom(2'b0), .bottom_right(2'b0), .init(2'b10), .state({trees[2492], lumberyards[2492]}));
acre acre_49_43 (.clk(clk), .en(en), .top_left({trees[2442], lumberyards[2442]}), .top({trees[2443], lumberyards[2443]}), .top_right({trees[2444], lumberyards[2444]}), .left({trees[2492], lumberyards[2492]}), .right({trees[2494], lumberyards[2494]}), .bottom_left(2'b0), .bottom(2'b0), .bottom_right(2'b0), .init(2'b00), .state({trees[2493], lumberyards[2493]}));
acre acre_49_44 (.clk(clk), .en(en), .top_left({trees[2443], lumberyards[2443]}), .top({trees[2444], lumberyards[2444]}), .top_right({trees[2445], lumberyards[2445]}), .left({trees[2493], lumberyards[2493]}), .right({trees[2495], lumberyards[2495]}), .bottom_left(2'b0), .bottom(2'b0), .bottom_right(2'b0), .init(2'b00), .state({trees[2494], lumberyards[2494]}));
acre acre_49_45 (.clk(clk), .en(en), .top_left({trees[2444], lumberyards[2444]}), .top({trees[2445], lumberyards[2445]}), .top_right({trees[2446], lumberyards[2446]}), .left({trees[2494], lumberyards[2494]}), .right({trees[2496], lumberyards[2496]}), .bottom_left(2'b0), .bottom(2'b0), .bottom_right(2'b0), .init(2'b00), .state({trees[2495], lumberyards[2495]}));
acre acre_49_46 (.clk(clk), .en(en), .top_left({trees[2445], lumberyards[2445]}), .top({trees[2446], lumberyards[2446]}), .top_right({trees[2447], lumberyards[2447]}), .left({trees[2495], lumberyards[2495]}), .right({trees[2497], lumberyards[2497]}), .bottom_left(2'b0), .bottom(2'b0), .bottom_right(2'b0), .init(2'b00), .state({trees[2496], lumberyards[2496]}));
acre acre_49_47 (.clk(clk), .en(en), .top_left({trees[2446], lumberyards[2446]}), .top({trees[2447], lumberyards[2447]}), .top_right({trees[2448], lumberyards[2448]}), .left({trees[2496], lumberyards[2496]}), .right({trees[2498], lumberyards[2498]}), .bottom_left(2'b0), .bottom(2'b0), .bottom_right(2'b0), .init(2'b00), .state({trees[2497], lumberyards[2497]}));
acre acre_49_48 (.clk(clk), .en(en), .top_left({trees[2447], lumberyards[2447]}), .top({trees[2448], lumberyards[2448]}), .top_right({trees[2449], lumberyards[2449]}), .left({trees[2497], lumberyards[2497]}), .right({trees[2499], lumberyards[2499]}), .bottom_left(2'b0), .bottom(2'b0), .bottom_right(2'b0), .init(2'b00), .state({trees[2498], lumberyards[2498]}));
acre acre_49_49 (.clk(clk), .en(en), .top_left({trees[2448], lumberyards[2448]}), .top({trees[2449], lumberyards[2449]}), .top_right(2'b0), .left({trees[2498], lumberyards[2498]}), .right(2'b0), .bottom_left(2'b0), .bottom(2'b0), .bottom_right(2'b0), .init(2'b00), .state({trees[2499], lumberyards[2499]}));
endmodule
